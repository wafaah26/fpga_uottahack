`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
s+wgaV8JVJYBrLFnk27HNpS/tBrJmogxdlGySSKoGaFeLvUoVY9WJSoVInXa56JEyfDBs2vMlRiU
FtZMZKz5qQ1uufumAlFoWvGxY1tE1eFwLeTxm2OWWL9tY+tuwSG7hpBEJDDA/BhlV99WTm0z2GJ6
U6MgTWJMtrB9sRA+lYJnF4PmEM2Y+a1dOyVsuJRJLHhMqmkJej09iZkvW9m97gbepid5A7C7UIbn
5RoxvZugkX8s0yqbdzMMbvC4dL9UCmLF3QebV729L+5xU3+eIeLAaaVSpG5IsxM0eAvAFqzPvDXK
tTTuQjNOGoN94ViIHKEBjsUvgLE/PNLjPJjVxQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="f0VVHKDiTBi4ulppSx9L4daeSbsSdXYQAdFWLIbTQDE="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4224)
`pragma protect data_block
JDgqM1tdI0esP6aRkYPMeW1yAJS+MBbeh9xoNS81FRWK7MWU0CFFh9pjbxguJIKxOGIF/r52wF08
XlalTMR409FN8/p6pLE/Hxo1ZmsW/lSVp+ahRbLcyE6OeUl52A4Dkjrc1PKWyJiB6yIcJ/GsxkU9
74IUdym3zi+7lIiuqH6h1DYzSpMMJjfADyJjV7DvbJUEQotOSmb5xQOD7t6dPKrZjuWpmTw5sm5f
MPsEewH0joivlj4wsbGUFHe+RDzmCOWgRqiSvVMvLCCe3okpq44Gomw/DlQVZdvTkmasYtWPFAry
wVec5WUFsCtM8c2WdT52wUiiyRT/UCt3BF0DCMMWl8YdkGPk4u95k3R0N5BVkgbnJos3aUrfYZnW
MwobCrOeIXpnLYr3N2duRFOLzJukIDccooX5J6mDmfdHRRiTmlXmkWbK1+b6BooP8YgXgYoRg6vW
rKOWhToOwK/C4S8Ef7Ss/+UF1ObNNVl6FxTiNx1lGK5Gx9l6I6OBBrFlsr2KlifZvNUOUIeFLyy3
y/TqpuuDBZ1QuFI8o+43y6VCkFYFOwpaZX9aLb9P1816XrhDVsq/1UCHrR4OTnEWSZfFbk8jRxPA
dN+K5z0qelXfCkyEOjp7hwChbMqHVjGu+YdV6fhUAlBcqiaXhziCAN0PgQRfe2XcyWkLg0mBVP2x
PD86ssshNYbGqpqScE4dcKjk5/uGe47WoLXBHXmmJ7jTRefjmKItd336xinrSzFp9IqoWGw07BLB
J/830zwkwm6JV3Z1n/LMoO45g1QmUp0Q4pj/ZKy2ZtIzB8O3l3+gSJTlPQiq/I0dEQg/nQ+CIgVL
+j2R94z4dBNJfYyUDjZWsVY2zmEijbue0T29R88eF1qd6JEewjOCPgDKyKBxrZT2acfAf0elmjqJ
v+A1aA4qSnrfQADU/tBmewLg4U5PofEsrESW7iBWvhYXUKf7EUrGfDwOmFOwdp/M8psWvWEwiQ40
3ek23DodqG80EZKtgpUKYQ9i+/6LujImuv94nZ2Mnxgw2GyAy/heIFTayXx96DH31yBPFtxOMN+6
SKJyFLBmiydguLyMA+Ly1fo0YUyBul9FkuKpz6EuVJB09s2vtEYlcEMY7B5UF/kQmqT1N6gvk+cS
IGBM1Aq3CkEuxf+LhhCBm8jHfDxxVvVvYEF7+dnKFn67y8YJ02+eY75HweNRTO60NewdUnTQVbB3
Gwdaj4EtoRd2gbOMLxCXxvFrVYk/xfpMHu5RwD3Xa6MYHdzgw5CkO/l3qdgwq7zwFyhd+UoPEVVi
0ItYZcxENNB3IR1HyZDjoTB09v/yfy9RPvS6gHrq5R8zTuLTK6n5UXJOtNCh4SUx39cWX+Co0IAt
EmWTmW73SSbB2zrCbagt2pswa7u3Yhdfec8XqW5FxvDgp/S2vs7I4losnJDHQV8ohOhcuIwss/by
EFyZDt3JxxQ0sB4XUsP/p58hIQ2RC0Ur5oHLFDOeLKh3qiu7XVU52dZi70vOD+t8L1i8a96AcV0L
SIS2x1/uID+u3MvE5JX4DTfyCE2I/XGnMJhLXbKWtOU6/OdLVLZU/2MUU8Xw316lEHCbceap+oEz
J937vKamuchPZPJ462ZzPklk8kL+4ZetowhJe4sPT96ebzrZg2cNqCFrXWGbcqzZV+iip0d7jnPw
nfJNGbd8h0XlU7JvBQIvvKtDI9/u+ELqADtwwA0j+/T1Lm8wReMSEEAvsEL5uTwU+jt9TI4d8IPr
4DJEAkF9x8hQ3c173oZU0o38cRfQ318cBDaMY3/JP8n4RsyIxSQPcE5Eswz2/3Cj8HuHSRL/EPvX
BpD6eA1bNJ/9/zccMop02CsxQVWXbqjnpO42NHyqclXdBG1BOqa98pAIdAtUmO7kAtEum0KgXBiR
gPtpR6SJG675D8Ru/4lDBjypB0rdBSMpVluhLMhm8QFmVuH1K3PFIaZeElYq0zgWSbn04DWstPS0
BOuwWYZuwR/09bPVmvRwTnLssC8g7l7mpOwHT4j4MBZwbvF1tqSJ+LJBwB4NpQH1hy4Lx1N3Xev7
1Umu2uoeOQotysUJVFHUuUHm0Bzodae27NjHCm4sy8+nzALZK/sQ+3zuZuuxCqgtmoaP7xz4kasx
66Dt8PJl8F7BuwjxDFv1PpYgfOOtRpiZqgkaij+pTvmuU/bKKDxxB6WwqxLYSa25S7yzsmdYVepB
OFf44otwUIJiymX+p+0QEkmnKbYI3751go/eDTh5aTtzsLblpCdYu/4ZSCSoZttfkr6fgcl8h9+f
S0+7zqJEfkqqtiiSBTnrbdrh87/pTBh8LhFnDSZd+VEjCpIYw7gggI9+TBK42UHLJ2WDVXd30eS+
P9Id9INB3BGhA/1dwahumD7TX1nwxlgNJ884A6pSXHCZWG7AMDdxrinpG3iWQ6UFu+vGmlb0xSfM
YhmtV8oBTemoluDZ34kvNFSuvHeZviB97Yg2swv++Dg2zoOu8pnkGkfKG7ygzwmtCDZUNJfi570w
D+B/eRfwcdP7FNm2S8EjbHMQnbbizYjYf83lCPTLcRAc4m3xUtUh3O69GSBBBB553l9DdJUekrLI
PuMiAS45UwuhwW212q9mC6tP+aXD4OHzI/eydFCvYuDAaEAPW+IAJlWGSj0nx49+gCLX2t1LAJME
kc+TsE3npvbATHuyxNF20/D8w1o2spBbUL+P7z+97uQ3l62IgV3ADhnRh3L3w5mREt3KUquTzzop
XN8bCeUbQAbqaVGIC8KoA8IZntY84aA8p9Q0tRVDAEvJg+0Eh5oJdejgLRmCXv9xkN8RvfjKHB5f
hB5dqGpz1c/kWJCuSlor4YMFtEC7Llg7+c9RmGOSsPYqyPueeAr2l5CLVomVf6/Hk6pRYU2joWPm
b/as3bnG24JFCeZr7k7nFIa30QkZVu9RmIe7oIR4b9EzKFg6/WKmHsxXxYlcCBHNhhwHjYxtqx22
+hh9zMwaoGRh2WuJzruFgklFmq01YpNdncnxf+7lZz7CL2cP7HokWpqU6RxP5CV553k7nBzET4HO
NiPVm9cjaJjuypj8uhLen3qFKjwRo8l2ZqbrxVeC3puXHpPqLfhi0/m964PafAndrlK+JT+tvSpT
W6nvXp2/yeewPK61HR+7TjJWpCobUJEXxlpOZ5yMf9L8RXkMnr794PAWTmGoN1L/32G/3b5guNzB
Y+XIYXuljlWO94owlTe5ZV/qPZx+hkujcGVsEPH9PkRLBJPuAMwNDlBrMaU0fXzgs3ZNyuoOTXWe
VA01r/KNY7YZvrpuWEtcwgGR/a8pckBzlhFMtUmB+j1TiOWWJK3s5lmhPnaXVJxVVyWnlqlUT4bx
txHCcH05ecnVg+OlJEyZWq1Ju8KMinW3Fs2evCm+S8YIqKtDxddVRpMrHlnzGMZixR0+rO0BS9GB
ThTaJW95bHA/yb9alDgvc/uUBPVIoWFZlB3PMWChQoTnFzzL+h8/GEsJHzyDIuridErAVR2tkdnH
sjdMG1XgqMOqjnlRmeXY8BHQP/655eyGtXn/fLfttuZsE9bc2+s7Gi1/4b8WbWAYpGK0+O+H/URh
A3b8ZJQackk8GBxCb07UlY1zxilzPhpVv1miP/3RaEXoYsjtpzexW78eAbn04YXf8ylyx4HxQq2h
AAM8VGX7h0CYXmkRTuK2tOeCD+1r2IxmeDhxJk+38Ka+aEaL8msTqVX9p0WJ/DR9W+dzcirFl5TN
iGBJN79HMDFAfMtXsL71okwXJE4JGCaBJLlzqg6C6r585V2ZdKTKw9o/2cdp60h9EMQ6E5LP7Jsi
yBs6IGhALPCTAGN2D43rCPTArOLKzvV2b7kZa3+ysVTezhsPACFMWw9zxP1vxKV8hAMLNS/Va5Tl
5S+PDZmM4Yifylz6FLHT71CMXLkex1u7zn4zQOGFQdTDZE5w5er7v/YAhvq8AhMWG9oxkY2ALo6p
L19zT41jBQ8MBzN8FFNFM1S3cc8qpRFiDjoFWnrgyL3Pvh0FlVOkw+A890o0G9XfB4mcgAatGATa
/unqOINS/VldADHRsQxZs/KGdSTGtLNIo39lFxfakm37xIVQEAgS0GbWCzYDT/8ObyAQtRH9kHAg
2+OSQFN0PKkbbbVw8JkZ84+AfICUGUfqDPENxt154PbtcQE874RZKgNtzT6A9Vdglf7Th7W8VO5x
rnES+s+IkTpEY693qr55yTNs5oz7ZVIFJdr+BF9zKDjHU3NbTPtrhKl/NjYI7rkB20PTwPFTsNC2
GeqscOtATRtGtOc6XBN9VTZvWkRff4lClPz0MC1DMm70a1j8ru+K8wNC/p2HC+lS9Py1k7lLPZy8
zDZboxSHpHX9b0x/OGGOwjdCtel4GL4FXwKUsbbcGrarjz4jQo+C4SQ2SAOs6A5MSZZ0GeF2Q0jU
GjlYNqjelveY0AAIfDInfg5mFCymPtGuJbsPtkFSBvJVDnvcNHj+lt6DTLoE/LBcseFtKscXs71l
y3W6ZGluv+U927ttunXhBNMjHqS26NPxyovWMko8uZs6Bq6Vu0K6D0c77kouf6U34ZKAO3VtwOGN
du9WxzXp0MieTQdp7nAj1qzx77K/pSWQkLNOSmxO11NCbMD1o0A0M502gZZhL/OvT6KRoNNPoXFF
TllFerzdaUx+IBnluvqtiACnUp1vE7Py9I/z/jkePgwM3XXXbEChureiT3Fqtgxkl0NsZpnsX7UD
rzbuXAFDXzers/FMPgjXABYFnel4/hiIe7mIGUuDjGye050PIp5ipT2oQr+S7DzKF7BTnNk3Xr9e
d3Gxh8vPJQDPsz7Dw6hCA2TV/vjkik+VMMaBRlVvQw5HILglJ20rSKMBiYK4MGDU20/id31PkHpy
gloaNhwtjpvCNE6QPu89tFo/lDql317rFXYkFUT4D4A98GZccX9V4iPodWAhW3dO+yAy+rjEiWai
LVT6eT3EDR5dPix1NVok4tG1yu43a1SNIJdjIJ3Yu9c349AZ53IKmhs4rr5TD9NNYqY/4X6u6QpO
XOtb119hVaWzxODlZ3Qbss5d4r3PsTp4ochR3tO0tN9knAT3O+NhUNJepyvI1OrLrvjvHK4/Jf4R
lehWkefopyrRGrCu9CWnuC8aBVt1FuOnnKbVwWu2yiVs6GeQFYl6igVHCjRqWhOyPI06gXJ1a+P2
Kk5GexCt7T9+KGaHqW6p3HaU1YqRzhiXmNad1bmfS/h6toYmOZrMvXNVNq1Annnvp2enZoUq2sEZ
gp/jzH17cUVfnsdkP780/AtcRX7iysZgnjWJA+oUy9IDqN9WUYsHDECeyjLJPRtGU9yigCuYoHFC
ZNFnT51/FxSw0/Q2t+XIYDV5vLrPXs1q6YzWCxYY8pTmmY5Kute3euscl5ji7MSjnJ1H+1+IhGI+
/Rdjyw63LIRgB1xH1rPe/A9HqjhAqUJPZWs5rejcA8WAq909AUFWRj4E3iaXFBOtxc/Mvzt7qRvj
RHlJnh5HZhFYIbJBMmudKdfW2FH465U/h9D1C29MDGJzaz0iDPyXKX4AiXMLElTiccnxWRDGDJ3P
EMekCiNAHUF5DdVzH4p/srHXPuamZ+yZtyjiXHGmPULqXaVAF041gdDw2CQC7P2Ur/eBTo6AI3ir
0xSoCTvk
`pragma protect end_protected
