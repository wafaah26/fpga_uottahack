`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
eoqc8nRUAy0Z6pMX+bk9X1BrfSpbAOLHkpIFgOTFzdAynnONUZivQ+rRN7W9YJMGejSI9ApCVlev
HlA+jn8WkYe5rhgBrWe2FScm+7k6H7jaJhz034WQAxblTwj/oaW11jEj184FL165d7ydtuhK5O5G
GgkTu9vjO3RBJaC1XWLSQO5t1oCMRS3tq0BuDryfBlHm05OiT+TuhTexYXM0uMjfXnFxjz+LLdcU
LCJpKAUXvJv2I8vMaeTX0+BeMicI6w64Vm9qlMp83PVma94eqdqoQriMdBsrJm5A5ZfGgABFJkrx
p8CRUFXa5ECNM6D2+WuFFttsWTkPZ/qeqETONw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="l0780hf8rPcnMQjTQtoRUDstuc9cgac90nT0WqHiZA0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2544)
`pragma protect data_block
obqBOhIA3JfTG6gSMtWRABwvyG6eI1yNj5qF4pQKA748i4hjuvm7jDOPTyf+SXDQ/W8CDz03QNHq
annd5a0J7asVkOiJNzr4TUJNyqe6XWjmP8GCLqOOVRO5lJIbr8INEy9zpUQpDTGFo1dNlemThenh
JhdHmOTg0GAc7n1YfdDn0H9/0vAQ5ACvtEHHhSS4dqK/gVe/nJ+6zH4fKGcXDus187A97MQxH/uM
/1HnW6zqfZKHEG32zLdSQJX4t9+kf5PmePV32LaZDGMPYIdwIekoUmGiS4tiTc388FVqS1WtCnrK
HbaQu8F3IQtOQsYBA+K9M5dvZ3NrlXG6Ogz2DJiMsvoaljF6qOi6lwl1Tkn/S63XZHtRUS7oSUQi
1DXljhMynlf836zvSyAlj3Sd0kNFRTq/eZBAWGhbCTSNm9oASY+IEyRN66U1AftY22f7xX2irpGb
AYlhttzFig4HUlbgiW16iPtN6bnzwBYtePJHWPh7JyOSz5tM+ItG9h4vDiPMXuR1ChsiwnElX16f
unNK63o7f3XLHRrohE4Nw5eCi9L2Jdjbsi21gnIkQp/S3+PiVQE10FWoSYDrhapvRBB1ZtC6yq8q
XebWZ5GQ6lCeGeY52KkJOogorXSXByElBV3vCwCmvHORv+Pv2GZxZanQ/DasfbYn0wpdgs60QW4f
gcJlv2hO2osunSmoX40Pth2OaaPuvKChd+tuWi9I9gHhEsFP9XjxWQO8AGCpdc3PqdK1vKc+h3cR
FXxCtZTRdaP709JZ5Co/9nFqhCXlBI0/54augYUyySYmRtEI7Xj1PxlueWq/wDPqfbKPr2MvSoKp
CjgtqUnBE1/mvqphj4p/Ysim0o2ev/1bghi29P84NYgHeSXEntTUzDCm6vEbUr1kk1XfijEsmktP
oXzMrVlgaNq3pZ5oYqF9hFVY3ocwyylDPzgEBFmzOsm3E89MjESDV37rMRuGObmAvvLR10OkufNf
frPH7vQuGLIAIZyBK20oVS/co2MMumMGLmWX1kVOW0HME8iaOEFs+3OzIuyGLZdGMg8k27o0NMGt
jkgNPwZR4I0OuDlBg0wVEAnLS2xfoIlAbYV+UryLl6+2pCDnEulSDKLn5kyyu2WMiIW2B8jfsCgI
YqVWTuFWMNohmJGaN73f73AnMj1Btjdc9jW1G2dw3YZ00zOBVLLgqsr3z2yaOnISx12TUWqfyw2/
OrDGu2s8sYmNWam3jYzttTIK6CPh/7xe7VS438Bkqz42b1a0GgneNdMJp8zLCgLLXf5BZzR5bjww
5mkY+Gg18Pxq2BpKxFcPsIgHqVTOL5sF9LUP7lOcNGIawcveiINrV0Qi+NkrzG9/KUgfoa/WOLUK
iW+LRtha0QIDhdpJN0SCFrIyzQ9IUWWZB1WVNcyUKWGvxgZ2WDYEHmhYmGsLz69CsfqgzIdkZ/Og
6/omJjAnnTgdSYqm/IhirImG+7n03H5qElw0H9eYaXfMrtiN/junhJy6WM/Z5l/WkbbSE6Z75qBf
kgdx+FGQkxPYYUrl6z0IGpJwhHtnNJABNW6yepwL7pgQVIEDgXrsbRTT+1zJyuWsDTzrsSbi/sE2
GN/HZFP19Oc5EU04tljQQOQH3QpMSCjyAFmdwwEheQqYdicaRF8Mzt2XMAULBlHsW/1pvdTwdC6W
SGxHsFQGudO3qO2p1l+cxnjSrDKOvr09UNmm7YxBmGnIGkGJJdQkLpmw0YbYv5MvrLjN+QwxpbnA
/ejH/AMviv85luHW2X+e8FrwlhjFqrI59bRSyiMW+hUcqckHmSnrPgpEXNzk9JyUfFVbTDUtsOlx
huLgGiONRwmpjNlQHzwYY3p8dFIdQ13ymGF+ZU2DTEmitHyCDqBHgatTgr7D7aydydwtM+qMGCNb
7o7IzoBN5mx3HxjbdrNafDJKx9VSZ/t9Cujnj27YctXK8INrwk0WWCKqQlM+Lkavco88ttGWU3kO
ZxHP6IU4Da74tD7beJbJNASNQUm/EqKjh4LyPn8k8TeMZEJI8mWNbAWT6Dx5iltyeBqgce9nKbPm
tWJZMBGcJ5L5iFl8YIfvogkMVutxFPUGIBiQdDQ8sM8bBsSfnvwaZowNdqpBzEGOAjUx3njSdjRh
QPgXlBPN5u6vJPS/N7kqBGU8Rosmrp0eYHu5oIQhbSOnpoUhNNJQusZYPO0/9xkLvwPssx6JTtNv
kqpqF8Cw2bpIp+VdYIHEiRBOKAKtTARZgCwJfgFuQ3lSi980mZ8XJyTBE9LYBk/8ZUmwNgQba9D2
afWd/EkH0FAjZW9Wtxyt1SIUTpwJfAU9ybgsnypQr7oIc3q4dGDdwZOd8Kim/n8NxwoU0y1dRXgp
pFpyXANoWd8pyn2jOjC3LV01tjSOrAEHUt+frSPw1VOLByIQ6IBZlw/S08MH3I8JspmTKIuj4bjR
aqGYAbcfTdurfpZKmIUa/JJ5Sr+gLEnYiM1jKeOhebbSuSGn+rYJwnSVXBHsOMOa8VUJyCYBm08a
tfK5qNVKfY4zJVLC1cpFWP4zTpZrGuJXISjFsX1SIyT2HRzX2IB9ME9U+BTEZJJk5iLflExNnTwo
/SX10UCk0eYRVzU9b7gQZMjdBzDIRIySMB44hstWX0ETKaLHu67eafoGZmMzPwEyua2KSj5PYRf7
cCo50TkQ+8vOIj5JNhf7+QD3Facv5sWXqCYh9xj/eTO0KX31DcnrmK3gSokhVrI1DEBn9LeI9Ipt
TA8zYyMcJ4ND3DWJRCeaKUW2882ctClu714jQ30H3zFP+xZtxMxxmfL4kATXGrBWxpKkdL5V9I0U
/ul6SizYs9nKMxLtal/auS88Qk5npsPNR+QkG8xraNfbECPsOauPL45LlAr3dSKmw+mMuAOusl3s
yx5MuTAN4oP5Xd+i6kIEbLde02pNYl8yFjYND7WtG/bLSrDeCHbVRRjcH5Bdcmxm7KjZ1DDr4xLs
4zYlYAFRBuC0wyf1o3cOcccAaJz5wquiB3Kn8UViuZCWltDPeXXT/LkDz1p98Nbiz8WRqIraFQCv
fipSwFs0iEaNDEnqSdZwVomGzsj9rVbJ2OxN5ayse7cis4gyiNfFwLEd93QdSH5K99oLOa1Fzfy1
m8C3+H4uc05stBavl5xaatemZ64lO5zKRkUT9/Ctap+WuKUyOwOIEJo2Zt6xmUT6ycOxY5Yy8I+S
sbNeOpK7FAqZmzuJ7jeR0ph2hli5JMi1bPwFuAdnHYYo2O8tDlBHDoihG8PcbuoOjtJNkQQZj6c8
AFghDUmkJ2n54WagnA5NtnbWURhzeFJFa8Aek4ZhoH0TI9up6zF/+AfG9uZtP1376WW4c3aYsxVJ
jERXiIVNjrBxWepEOVFSy8GAHb+N3qr2XWD9uzxxir1YXpE+
`pragma protect end_protected
