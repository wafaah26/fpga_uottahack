`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
TN3QnZVzFXgVSePjyh9Hbg325HWDi4GNRngfLMoYK0PCQJua6zNcg/WgG3+SHWr+LfPq7jvysh6G
c2G9okJ2VeBpj7fgdAuzWfgzUnfuTFaqb53+CT19ah89rVm3DA6wTtQXdnMJ+6mlfSZul+DHlQwd
axNgOCoRPsOb8637T2VxeuZWe1zl3PN2rfXEJ5/wTM9st7sDdAZEw+ebGJOVt38naXWJ0JtUjxte
FOGORNDXtS3WenYfThfKddKBxHyeLgH1lomhs30VDt3Qx6JVBJvsd3jt+C252P+9ZsE4kpb2mFv5
Of2l7gRpywRtQSwGtGPV+PUM4pxaELH7lxmPdA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="R44hP4C3guHiNiQi/2L5C0MuMh5H8HV8oXCfcOtfjVY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3648)
`pragma protect data_block
xWN95Wo0BYiJKrjRm71/p0CfmFNDFGcN0k2SdMJHmpeZQX6chUrOWyGMhB4837A1z7GAoDULPzan
kLBneae/BA+/w328perJSJzK74dwsbomPpIOY8LqxAP/uI/gxHPsPw+dWBkwzyMB3rfsh5EeGZdl
+trnuXPKR+EBL31P7eDaf3hKayyp0VBTGb/FRPHdKqjJtMCwcHJQ2eXNrXXKX++dA7/J+1rWJ7Iz
eFjEWfUHVnW+5+XOMSIm5tYvoK6VbuQroRxCXxSCjXogD70VDMEgEbDgVAWqYONmw1jjU/norS6u
NlJMvN4KCzcAgfBd9KC8StPIZ2HuONpRPV6E1nNO5LOD0kmb/JuzPwpX+hgPdTQlxVW+z/msFK82
M2uVHTUMD6Rd2VTjcPzB+Pxqph9pLwGj7nfWzkSfNHqDy75WCVIflS0xJveunDQko1is1TAVh6Wa
CV0CecyVGXy9qao3b0zrmdLDlGQVjnKtQrCZ0dc+uJvzzEHYWrc0JxotJpDxeB5gldoBGr7zYl0T
l+UlFfsSUGRHpph502IiFTHiMvR8oOuEFtxTRBOIQsxBmmOT5Ob7hbgQnK9I9vMfp+BF8qniG1np
tsUt+FcE5t7T0QHcwPTzrbqo8f1PZRHRyqxFT/IONQ7okR3euVtmaWWBMafV/RREcRmAybNiTB5a
OsIKiNLZbYtxa+/H2NNfKa6PQgc94NoatoZzE4Qr1F6fNvuDYigqVGZFHi8dz/hAW5uC4ZnURatJ
7NJwC9wGHq++gXpTnT7KqRzGpZJhYz0BSH8ZuOno/UI24doTEYqSs75MIwwPxYxKIxpAhK3ywFOK
Y4Qf8FAN0FogLPbG0V0QELDmqH/7wzKjqtTxQhPTNh5KihInjCZImWghYdMOFomWCRG1Lv7Ljqd8
7naq+mdFHHMzdPY8QJsFmFsfkjJ9c2+ZddxT0iESMwfzAZyJohEzy/Cb+jpsWMz9WX1NFpfNVPTc
u+kZomh3NkGHPsqAX6kc8F+QwoOuRtkBrm62q188IcRa5Ch0+saKpc8nxM3eyxJ+xzhL8a9Uub8L
pCbS5W/v3kfmcGf7W74aNOEaGOuc/m2cqLqTiWj9nDzeN6dekeQ6NKof29jmQ7ToYv681SoyeIkk
QQIas9M1snuV5aSaSoI3Wr0D3ZNtf6CuuzmbhnnVs9d5oviQ2bB/VxYkAS0iDRyWN4a7b2aRDUBx
FJ8wRePb5Su3/zRkpyNkAVwJPCRMMjlcZQSiOJAvBOHTdpMhvzYli2rUoM7HNYEAHeCZX1jB6U6d
bBrtt6v1ypTGqVeGQxG7rEzNXi75M3WI4o69zEykx0vMa4kreNCnKcxVDe/xuWhrpWE3JnjZCTMQ
rTwCI85v1fDb09XrYTzZm08m+mpjPmWN9Ao6o1utn9WDcCVWL0LefewDsDvHrZsO4PTeouR3SJrI
aW2zgP0tVZ0AVA+OcSeweYgpECM1AF57I+Fj68eC+kDvnBZPpHtD0MEwRzCfC+jUddutmqJHLeUV
PdczAE8Q/GA1KyZW4ibK/Lf6DuPdvmHG+caP1+I9NyXRwn9Qb5/ExUhjpzpB1S36RZo/Jxr82jQq
rBHrtxDBb+kc7rwCyDzVG2iJf4kcIE1YvJ0cGGMtge+scRtwLO/dd7E+5eVodaZMQRFKhfnNWrQx
luXBlkTf3PJdkfriX/zOeWzFcfH5tgTz2Iwol8qRZ3ChbDsqQ284yk4yCdrldVYZLdYBfCteUFT0
PIac8Qqcaatukn824j3EdqDfHuBVR1+4VzHcf7M85/hCCoeymFsnhO+Hw1PJCoseH1wtL73HBb5Q
tqczrjhDVnjnkfq9iF9zSHKRnmD0oFoKjTjovXtqq9qaowAXskmLP/DsTqa+I0nirywf8R0O3iCN
uvO3xZaJsRmUp9h9xX9Ag4aSQF3S6hNYAIlx6fQ7+WkeG2NcST+ICDJkd2R5dsXpHl2WGFRLYyIP
5vKSI43oGDF6SBQ1xJyzi70JP21TAr2Alr6WW66Bt7sSgxd9bwT7gCN5Iw5BwL0FJnB3u1eJW0N4
7uaYFhmKIQEsDgTK/8bOgVa7mr8xZVLXE/1loQ9Kffs8+e3DZ0S+lSkjAUFXklZRUhov512XIKPa
j/yHrxZSYCojvxs66WkiD4vXBT8dXFOQ18G4tmdtssG7DyhHx9JDJJtfGF8gVk67iOdDhn4Qj7sj
O8Q2yGNCF7Lmz2hXh037HUb7EL95gDxEGW3EsqPE6bMjmy28Pa8Jc5HCvGMWgItQztisuEI3meNI
88IHsDyo6ISu3SeOa5E1hlhXD489N06SlKQP2n4nwz1AV9Ur/CYRaMEkuZhNr1i0T1NDddon75pS
ZvusOuLUAbLShKrN+nsGquh4R/YIzj3YmCWh4C5ytUlgL/0khyJJi5Ccml8SzxscAGHObC1IU4vQ
/0QC+o37jcVOlWmjUzurmtdH16kSUIPivtN9unbHJZPIPcmTWwyolYagDsB3plxyyc7i+nqO6qJ2
mf6ri6m0ic41sOtU6XnjhrPcgX5f/iK49xLTTSNApaKgTg1wyusSy+6rNBsTPez9aXmlRaoCgD/5
MccXKWWGeUsPREZ8s25XjmGe109MdkTrHQf8L2NJ8iwHKoRy/ETCTWWELTKd3z5mH3cK/OOsx9eK
Jnxh/ZKL4mXAKfgqjYf66yezRIRee8G6ccAg53SI+Y/NJ7mKV1rPfQpzQt2E71q2Ub6p1kcD6rpg
CfsJCxELWVuNaxX352M5o4COfYaILc8KCl/+LXlXuU/AvuSQM8DZZO+8xoI2ems75hNsF2pKDfmd
HXZsufXcX75oyWEdyp0RpKUOj8HqGOlFiwQKgE/vMsIXXCXiHNkL2bU2i2TiaTStg5favPbmtYaF
FImpnQIZKiAMBWPvQ2gvXzT/5Sx4gnhZfb/NR7DE7dx7VHofD+u19KDS74uvdTC5Nk9yLQt3mbnG
VSwctjJjn40gutcLFoLuKogzDTU8c2z8AKsrDo4BkklrR2+oAO8sCvJXZGaJLdfYAF9pYxDCCysS
Rk3ohCT7KEtUgzz/cnNjzWU3bObOvCqPhZiIFb0h5toAXcRZzXGSVLeCXK9keOVk4eoTXv85zyWp
cvJiKcrrfPoxoZRB6KAgcnHVwLEjEiJSmoqDKDN6y21VmEVhFuad4w0L8VcwvZaBLyIf2OL2agIQ
FZ9jYMwXZle/aVM7ctYon4GpLmTPHEPk4rByBTxLydmcNYr5WASLVMRaAul6HGDcOpQO4LBqL5vq
ZGzkG6rrDHiBK9aFvRE4FQWv6ajSgC7wbLUD/jCW1FGRubqDmQVOYgd2H2ej+xjKTc3JFppt4BJ7
9+kjuQxDwewMZAveT1olOP20y8EpitQc6x7qlaVoULKH1lJdUbPq5PYVaJePsILAaEmvZiRfVEGT
HA1P1qnrjbC0qT7WreOSzjuk6xXeOiqe1j2GTrAEUCQGwsTOQlhVMDMtWHJ8Clb395xm3lFpZNA1
1c0+8HBOlHFbyBnQKvfXc8fN0u/970245gg7QQNe0GB0j62BSDEZA4zAc5wotINRRwOMZeKHYOUw
LiEhW5O/Y4/j5o95QZVVHdGOF1Mt0LhpA3wUdZHwdP93CxE6YY90tW9aZ019w0FCgmzsQq4YM0+A
ASnGjGhExFQnJDp+D8sJp1tfxhDZTjygV4SLWSaKKFfBTxX4RIcFdY/u6WJcmw/iAXZO6IfMf26w
M/BJCElCrgdPZ+lk1fA+clhI8hcSzZRkGCRLx8Cr3KFVhwvtc3NFYSeZVTfrCvm8jMTQ7RAgmELg
g65QBXXhGQlf8YzS4+hi68pnkIpLRmUn/E4h9QczgjiwP2ab6tfkK+t/hBvAzvSpclrd5EQb94+7
5fP3v42fWWIcysCEtZ2gq6yFR4jaUht/8SG1NpkBZBXtdgS21IEyQ0cbimG4CxJRyiflG4IdX5NM
L6pZ53c8Sxi1fcoszVuRB6LGAkhSEVJvVtxj+HacCSro1d4G0ZxHqu1VcuaegvVHT1lc44woDBlJ
ZGxeSi+recYX9Brz0+am1iLQBaUF4cROPyhpaItnQLEsfMFB8ig6EJtB6pc012zv9K3Gmt2sjSmQ
SHoU0S4oa95zBxXrOqXVT4sIgqYD1zLQmZss3qom3BHq8xSbSP2wIwigbYtNTbuu9CgLmZCZVeBJ
nLk0EX81QYQMf+KgY39WghvK5ryMeDAKxUv5J9+9ok7rs1LWboHBmDVQUGTzECWvTHUaSSRlsNpw
yDANlH1mIGdKMty8d1vI7LU3OEbTIYnOkKEgqEcYG3/7+uWJ26p0maUumyPf+tLZ0ShYZRRt2ApM
dxv0ytkyOVceUK9L+m7/gAvBuOoyAO65DzuLh8hmuBf1vjfimWQBnnaOUqzgMGljOFgDNaz/izDa
JIv9gpPAwlvboQ0TDJ8UGnXlxGhGL4NcGhbZ52Vg983iE25VM2QKtEIomTK223gbaV7kZFQyYoZc
2laKQJBnY3CuH11MBUtSXzp3+auE70shXAZ/N0DrpRnTD/0vsM0HWyW9SAZ2b8MCprhjpb4DF3s5
5klKvnIrXeAH/nJkGW9mZDrw56WgylMd/KEl7O4bt2VTD8VnBklDLkp6x2xZqDf6CFNoIT/2BhNR
vqwdo1mZYBCGOfJsSvjrENCrDJHH88TZegi0gO/gWriH834K2Yl+iFXXz9HW/7VzPEm8YSOZHnVJ
oZll6MRbEptDOpZqf95hAlPA5i8BD8uYoyok/Kj09eZvIBHmGWNEEpwEmtoFXyGeN16WsDPMs8JR
ligpwUPSs37wJjsGJYCPFn7dSDUXDjEGwuAoWlUqrG5XkgIXS9FX/JWxZKsh+XZlmGoa3VSopohj
`pragma protect end_protected
