`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
dXK568Ag5khg5pdTbVnnYf328ab2lnTpyUj6pqRYGxO1el9o6ri4XS4yZNv7brZY60l8HO6EVVMt
8F8kGNssOhpIGFXv3k8yZ1mBxsdesXPoHfyx1VfWXvyOmOiMk8NkerarVhJAhg6aUCd328lunAr/
LnnxY3QDRYwNk5aqBJGICKgQf3SXssN9zg7O4ZG2NOg4ROOuj9OB+BIas2R/U+Gn5XefhuRTFpSA
n5uB+xDtEGLuFeA7ypR0onXW4YTq7Mm9UuDyuB5dGPoUfx59kbFx1br5S+GdP3e3FWnXLVb/bYHa
z5RP6k9ZLg5ZjjUy3ld0eM7i24WTgrTZ9wpnWg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="x7dY1OwrXmD6UQjYbQR59ntUaQrgEFPXmGPSon211k4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4976)
`pragma protect data_block
maDW0wf9IGTu+M7kkKyT3LjuHGrVYIfiAEywDjg1DDCBMXBCnuIXxf7kFEMvrY6DgeazRYkhh1/X
8Fmn45egEoL9LPH8z2gFAnC3HmhNw2pgJNeuvvHHdjdc0TS/BfSVdQbYApj9B/da98p+2KgL9M/b
bAwbEWBT8nReWD+4oxmlXC73EB6zuRLyBF40wMYYAi96c9HIEU1t8qPG4EsFcaZkGWSDTenxPPdT
k30fWoP6DDi0Ye46mJx68y1+f++K/Wp6UpxyMtkj4Ee3MNQuO7ZFzabXWGbG17tutgAt7JtK0vmX
/veSwucC37wL2tdnCM13c8pJP60jJ626GPXzB5BD0NSBR2BQwvVH2znqJIM8P4faH5AfueJ2dvaj
JeemTlIEa+yG9E8fkX+4O1/AYuWnT4Dj3pSJuczdOYO+WblCsyXsteKNU1EVOMLOLBHPOFSoAQFV
vS0U63RzXHYMO/IQC7XAjWeyFRvrcxPYlXDBDg0Q5XTVy3o0Fo+2AfiCFquw6B0kpX+//fqDSZ4W
XBvf0HVQ+B74IE8McIT/xxmoRMO0B0KpqpXyAOWkIVwVW67yW5TGtMnfnZ4aoLTbK9iARbFAfDza
ZLUCEYCsl/BObKZWLORulJnc1ar+dk8umZhqVlW/FpLCKwZTOKM0qr9nVwEBII9Z6b6qFciUmHAi
e+8Nh7F5XPww/ok+zKbdZP+s7NohWTMT9ok3T0jLs4uhjewg2y3FUaFX/Ya3kGNFlNr4zqHF2NQY
G65igf1ufgcVXXgncTDD+pHVX7jvKSvMOQeZjgjJA63mC5diyy0PDuJOxqZ+slcfSU3b9U0y3N5k
vOe5kO6kHk9MvNzXZzCRQl1jq5bJcqKCHLuD6Cx1iQgFKVHWKXaBhH8EHSzhenB1MqLL1wsU5mOl
v2Qi3IhWei0V+megZ669OBTk0FLhzotlh0E7xFP7fHPxlIahqWJ5ussuYSs7cvcmogTuW+rrJara
MyQ5pUk5aonNcsYYwKP4JS09xARuGwje4uMJoOqcc7mKMAZjrzZR34LGso4fmQQcVYtSnKAAz6Oy
GqSibs/EUw055RiyREm9MF+B0PQl9fbghaNFnxWkkVg9pv24ppNByJ/gMHrndfETYmGU45Wct4lM
KCppy4lDljSSb4AJlc70KTfYz4Jw8ukUc+20+JK4tIQRd916nRoxj7CX01SBqjF27An51t8nPUhi
3VVH9eXybtRh2ccG9eFFveUSaC2z1gZl1grvHAFD0wLhfimwwU16PD7evCs9k7jwiVMGPp8A9BiM
9XtdQweUCtUHDA8qfYlpLWXWxp+UPlw2hPv0m1Iu/01r5nE9WfFtwUhvveHRw/jp89Y176TPd27j
jaA0JWq5Q7o7QKK0BW5Ki8JuHYXqZsg2C4suZzJslXpGVbFitKcYkP/EpMOdfY/ESHQCiHFDO1yM
OPR0ybCOfhWPAi3drn0OTKcj3Q3YcCFgMEwtgrg0Ej2z0aLSIiJFCYLd3DjHxCAm/5Ypw6L23CSh
KI3KhnwYxOeT9jCjSV/ari0sg3yvztKVgNw4UnehpnxDYI1Mhqg6X5nteG9dVi0SWbuaQ0WZ7090
nl72axte02mTm1iQesINirF3YouwJidEiLlgg3krrtJMdv0b8yHTUiGl264k7HFSnH1ch+VD3rER
3CLtxmegLHnb6VJoDfBw93t6j8Z9qwKhSZOIMz85z2we3VWFa+3D8GaYAY6xD3A5YizA5nYCDR58
Cx728TavjCND2pPDq0Uwa4sQRLkpMGRDM32K3ZEVUs3KJ7IT/FYw893RJ3dXkFQjhZMBXAO3lrfl
XDN/PhLkck/Ume7+cKtFGJ4BBAXt/TwVqPYljsRCf5WMcYEbHXt7p4vUl6EUFEre5FKC+CsIGT4I
ZOkO8RYHmI+rtu84BkN6zHB/Wxeenp1nQ2jjDfDIbSBISScx0F7l/leYYHL01jCVLT5+WLxTEfQK
u6bmXMDGw36mAdU/8rikdesKrR8HOvlipmA0TI9LUP9t9N5az6kJanctQWV5bQskahaZzuWy7lGV
9AoiFeMbxGRe0C+n+kUl9BnTGdOvSCFng3avOVtjjlC9ZBz6+ntsGhL9nE9Cy4hN1ZEzw4IZEOpz
x1yvXOn90rmp9hX70Uc/jFNM5jMqhaPxR6T70wQgKTRMBHg+a/U1KvOA8SmZWXEBe8rzZRcLHrqF
Ad+bAtHOC+V2NAb4XeqfJpypj4UlzZW8EITVn+3qz7hY5koGcwQpcACM/3dlsBeEK86sr7V5HJUJ
kTZAoiTrN4j8Jo7IQIjybEADGr4r9+MJIE2iYfRcOTbremcsXVqlmwr001VKHNAR76iqNBODWW1O
1Cva+Kv0PoGtpX3zzrrdbOu3km//8m6IhsXeF0fBVksDQbkwOS+m8erVMb/DG1HelROuTGmiXvzL
AM0GWnCNkd0JXT7KcwHMycQ63kmOMyEE6WcMbhh3ZH2OyLHZVwClGS7hvA9IeiVPOE0gNl/oLDGD
soJ3c9HyQmJVWXlLCu+i/TFJ+jNBIzZsXwnFnibnDb5XhK63EiNADkuy8Q3QTh3GHtJSFgrVKh8C
FbQLZ4Zmv7rQm0m8CCSG8hMulK6023QymaduZ4k2sbF/zruqDKP3HM/bXytVLo6PcU+F98SoiLAV
wcE+LNIyTD6MqqocEPbfDMotBFYG/J9udaMuRt9tdiFK0ybj+RQ+yQ5DiZMsluz47foUk4Hqq4et
QrIeCqiPGayZns5JkWslTxQymeIciy2VMgAgl0qTsoFwXSv/kh1+4vcUexTcj+92uXQKHwlUTgNm
inuh0x7uyDHEm6ABMNR9d5j9XhIfTfedav3CwPz1ACh8gP51cA3EDZ456jy+s/DBBY1CsjDWpJ8j
+2CHgpbEn0mPMoo55fra/bwnM9OUSRrNOZ6DQBpTJZNKSYy4SStfyQ22Vx+S1ro3mZdN0NUOK7JI
MldDtvI4fdpltL2GsruOMmMq+neH4WjrQ3Ng+CITPJ8lOlXveqlcF9/vSOMBKG7EsmzI1VtRVxuV
GzHTlfbP+R6Cz/JsLX504IlD8ZtazIodcefEXjs1z/ugA6UFcHDyxlsF6thFzh2pnAbt4qoAoCeL
To55B6yEqSuT22Pm9FEJzJj4umYHQxKp8yfOklcGFONWidwZm5ebzT4I2gKp5DZ1i73nJXW3nf/A
S7UauOK78h/t6z5gsZ13LZpxUKpuoZPw8xYa+5Y1ny6qxeKKlpXNt0fsKwwEPNzP0rRaRqV9SIZR
meR5rtmCCSt+qu9+jCDpNqKzD3sYUUnNGAcXp/FC/0GmByexzA0UTka+ArrmCURxlupOFff9d6aD
pcO/yaHPNm7hfybKq0NXsT1gplvy5pHvankhvSvLmxNeXNClsjlk1c7OPr80n9WaKeuADKCW+Qrk
ZX/xITkednkj7blx3EsF7/XtQ2O/74brmc5JNtchephZ2RdhkP2WIe+BR8a6TDUF36LQAR1KTzl6
2TNPB4I5yjqfJQWbjywWiC8m0DcBoJDECM2VejZ6CHDevToDPAs9DUvUO8v2L9wm2MLcW/CIp9Oh
p0JUHerE23NOSaZoUn+N0NglWL8X9Y+Nn+Pi3vME2jCOzmF5tF11GNCvDDXq444y5CehytFtou7D
wj9XvFJOec2/7VqyibTpVn7NrjFZcPO8zWyCN7++yEZT+4Wqc/cJKEjALH4zilgoyOsBMBvpyvaT
USgPBU6SA/OQ45PXZ3TOpsVvLaDwFxDavh09Bxg7mM13H//rZbQQ51QnJgJHnT254+LaSedfcIU9
XJnASFY+9WVpHGka95/9+3Pd6AC8XPrFPuV97JG03LOlydJxJq+VU4XmR5442pYXx7wA3sK0B5r/
3rnDOt3lFzItT2UyzPLsbOwsS5dfBG7SLwVKC/lltgOIumxUFYMtrVGiTDWDoO83hkvZ0EJ0ZlGm
PpM1B6ukx4QBP9GpBzD08vS+/pQBodNGkPN8qVXRAD0/zoP8wupL62zyyIUBEQz//JDIvy0IL/RZ
ZrADxp/lExS1PY/SZ2DpgZU6v1rnKz1wCusWBAIkuJ1JRKL+Rca/BsJBFn5OmKi8yvPDhoL4ktWD
2sCSOLBYadpjMtqBEVnGduSiqBEDNvIWepHqXX+DwMtWQt1lEDuzCtHiwOm1dL4rzT1d7UokLYW3
oR0udIe3eonuLgw6tpSSKQntSHhmmy9OssTUkY5IehHkKJHGMAdF6nLC30h+pM6eeiR3Mx09j4oR
hs/3FxpUcH6E6mUbclgkrwf5G9M++iBWaqw2rPeCNFNNkJCHh6WWR6s8DQ40STxHbRj+94zz88Rd
W5sOPnT1t7k8RoIcqYmd4iOP+jl2WdvC572fB7UrLT3uKTaZqcptspBqc1s0Faz1UJO+8qnLpAFG
uh49Hyp4U0NuHTfVG1ctNZqaO/gniswjyIKFJJxA/UTePbrKTqX/JquyRLAbz4U3HIVrebm1+8TX
U7tj8UYEC6hS8pK6fVV5TeWVsODOGvdgkLU7ZfrC2TBhKz2JG394JrsQS65FG2NDd4hxcIL9m/Bl
1QcWKqc1Jmvm5MMJEk1iZ7hn8u1k0QSMt/nQ/fMjk7rDZ4Nz90AsILOe7iwyRzhqSstV5vLsVmrI
UeNLqGDmWuunZKM4qBpwJhVQ1qVCbBiQXMwhEawE7wHsjHMV92JKRObQTdpZ44TJIq9Ax/Uuk/7F
kfk02BjlpFXzqERaOgzvXPbwaYEjYnx6oZk7jqdTe1ejRfrwfZ+3TirjLZPxtEh4MNpm3/imGSHF
pUw8HpszjRehgYFAfqNrq6M8/Exqtl6Uh4Y/MBKv0n9PHx1w/mJOcawJF111cC3EgxLsH6ot7un3
QeokwmL1NxNJ31cv170coWbWjm8HfQvFMWItJc79jFLlIGPCN4upjKEF8fK6FLTjDeLdkHwIwTeS
rASpILnWoV74OREKWGVI564jgsfoBIKQPZpUCo76eMxZKH2it+AQDeGXHBCYuDkf3pKH+Yn62hdo
0E6t1LbpmfGGz6rWoCqc1yCzDOCSLHQwJ+wOyEwuoFBZnteVP93JwwlqPM4sVXiRnPCcDy9iV9n/
vYSc7DyPac1LyrKY6SUlFUdz6E/p2uGrJsoLHzr/ABMlpKjvYDek0cm01xl/oP8X4+9NtVOqK4Pr
3LwWn6xCR1TMPk/yuG1ubjEQXN2gyxRgI98oDWuQp2K1R7U77nEFHYZh6NIjmILVyqR1vTfcKtJ3
SMObpDnLLnNnJzreiZoUhbkQ14x7jyxgqYXEkwnDGAbGCa3SJAF8aooWzU6LRhPNKU8BJvCyI3Iq
IKGDR8D/7yRzFj7Yx1OcCn4D9OwuO6XM2QNaRoJ7RXPe4UewY/R1WvRUXle6N+4xsSvchDPu+vj+
X3mx5KwxCCjlylb8vSQJR0DoqeGMJo0H5aVo+w6pkMs6SpW2GBBa7aoNSJhAvQsBN3TuZUcnwcNR
oQL9qgQwyzhrA75jjz/eO7YM7L1BMzBhuzWEJMmIValFB9tivsktWMro4XcV5quc/A5Ha9cWPFJ0
Sobd22lqfRdNWOUa+l3PV9YO1azpU3KoQvh1B5rRq8PMLdgzVwNgX4cmBrUylJGdOVY+yp9i/6wF
yr4czb6qtz3J6ycEiFD37+y2aeTMzxl5N9cLgDLYVci0nIGAbN+V9FGBb/G5fsabvPMJTvY7L3+w
kC50wKOqW+SdGPqiiTuToKAXHhDHQJr5GsEoybNfxk7a/a5m4xfXNZrzAhY2/6Eoioo838Mm/TGz
zYGFnC30MOWPQ/scOj9XKIOgZ1HbELmCGo0iUO9LC5pqAQuNFgBjA0Sqm6nRBPEuI1H5BSZoKHBv
a6iiO1L8xt9EdiSG7dt9OjcTRL2p+thRGQj+dau+toEaBWiUprocgSXOVUMDTk61W1pbRpAy47ws
y9chxGUl7QF97F8SPkvgq/oBkyG+GUg5MQtPC58ju4DnMGd/4fNICJnAQOUmIxUo9njHjOGGfsHF
JVnZDAeUfqqeOUHrauK4fuXnkxbF6oxMcEAt2SYmbKqXCpIebwJ+wBIN8EpV0F43VMrFV9wZuKFP
iOYzwVSsapyf6/tZ2x2mbxOxsJDxYzN95duCQtL1yUoNH/F1NwAkhvVTUWfpcpNtbBiRHM/KONDu
zyvw1FecC6s3VoMWrHe1RMh79BZwfv7KFEQPNwVqoRlt+rrmLNm+njpc+TX73E3oiPxzZRyRHWy5
i5diTyEMF+Zt0PanlK/Tb/SUhvVWYCdEUOyd2JJOP3uPvOxbQU3I7wD1g6yKy3lOgdGjS8IUdf8z
27pdw4HWKjwqPBtjTLxQ/FSJ2zBfVFy0AVIDYlEMnWzze5td2QK8Ioyxc6pz8AzRKesVY+iFxcsF
mjw8LcJBNxnfF86AXbr3HYXNa91VtpdHWkmtPSnMqfphELNAgFy/XfGHUvN3RqSySPbwXRkW0aOm
cInNjyDlaO7vr9D0HVHSvt99n77eeff9K4F6WqyJ54iWwMdZyQuMTq5RuCso7q4kzXumMs2+Kt1v
bpFWdaAyFbZOA81Lng4tjWtoX30qHCsNvVZpH5bi6LCx6/fLEs0fzlGPszNneaUi9/Dk2fmZ/pdA
3llzS0fFwVoTPOWui2uWlSo=
`pragma protect end_protected
