`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
jcnPBvMLr4mmY1qTRNY3KQ2Uw4YUyBCAWBaYn4Si4asZUeY6S7qvWB1sBY053IycM60zlusttrod
AgRKAbbaMzl3i2PxNVHyRI4SObxdm8B699t45KYyeVAECTQDTeescnYZqZB1Pd+yrPEz76/8qVVb
Mvav6mtnvU+mUfBXmcovcO6oKGQAYkIMVfDwadO0ClFab9bm9X7BZUXlSWt7zRcxTAA4L78Eb3uq
FJx5EWddFuUbLxumHGRLc3DCVo+PhWb37duYVxHGKlcoVbZA6fJ6wIAkydaMcrtmAc4mWMmYe/eZ
iSeR0llvySAoXx9Lxwf9VBej7QwPAhXkewORfQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="dc2PlmLEx7A3WZXb7YGdfSdhHm8E4g0Bk3IC4RRcyME="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4480)
`pragma protect data_block
C83e3fVjLUt7YHJ2XukCq/aOPpvD2ajtcWEf4bk5qLte5DNAXkaSuEXBOk4yz/LXeQXx9B5t/mAp
ipYWN7jJZ7Twj4zD04VE3dAHDn3r3SRhjq/gi2+eIqJr1xasQgM4wj34mqJz3DO0n/I6w6pm+Q7m
jgACDVMAUQJX4qCkF5OzgZyqiz82w4bcgqq8lkR1yge+N/+E9Odkh3BPWLBWBUwSzLyfC6AK8AnH
ya9iwuCOyD96A5GJgD3Vo62ElaHpKIEt8cT+LdTNP4WuFEOhIPZukuNGULm+CeGW59QwQq/N9S9t
H1TLCPGqcs3MRW3sFugT/6syqM+2cGYt2no9EVdAnD5TfWt0Vco/Ry1ULyJEPfi7L60sIxU4GgSl
dcJZxf66iaz8wBHXPTYDJ9Pqb5MFwiYSoq7h7fKAkVCOv/IQFBDNDU5NdnOqNB7Dlkn04HB5Twih
nf8TC5CLzyVytqjYiaCudQgLVZRy8x0ifncJ3s87zPXlEmYmZVqjkhmtFssDBKMcpGHV/SYJCu8/
vrqOsAW49I47W+djabnREcSZepn9DhGsicheVO9AMK4eYnp4FLxRIwETJS4QSV7jz/dz9Uu5ojX5
AL3kRr1YAUNVsUnaq/v2ZaasqcNqg8p52YjWOOjIm16iQmqePe/II6oqeqKaZCJGQit3BWfRHdEW
zHX6MXLaBOPYcDXg63CqqMUwtNVMJW5HOeoxXtL1kPN8QkceZ9+jmZXdjJ6vnsyv/W0XXs3MDov7
ddclQpHaAFvj7nQM2Cbc5tNm9K/4YTikhyUHgoykYOISFgfHSb9JV5CH5PVytbQSE62zyROaDnX4
gM7+enteKQOIDJA/b9QhMNwnRFwqw4crXDrydahphf/yDnBGGkNaEisd7azm1U/2+VpeL0ziRM5E
AyRr/FA7gY/kg9Qn3dadW3h6HBpbi5zW5XWhKVOkpqLroI15wlTH10vcbxducdoEC1H+JIdu7VZs
cYSkvvXXgUeGlb2cK1H0nuXV0sc2A7Dg5MhOG9+3u1gp6R1r2eJvCk/GJHuKZjOqDBXqXxdiprJ3
LZjk10Z7H0ePv8yzz0OEm+81g0M7q2e4/nyJMODWT92UKcfKerA17u7BwnXztQRW4kxti5cY36Y/
Vuh3uv3bem/t5ttjsMeGeiYMVddG4oc7FCNV7qDCMmYLR1tp+y7HTdn6r2Xebsr1CLU5rL6YjD6c
s4j+6SakAkqfMdY0XnPdE/beMi/zdoXELDQV6fnft6jRWIlWcUwPfBZq8FxovNC6C8gjI9NDH6Zh
ju5N/c20nwAZQ+igGIcoXp/F5jy3hbGYw37K6R4KT4r6W5uo8UVtwzYg11hUjfnRiT8q9O9qOfAw
cGvW5FJJZbeT70m+IRyRFw/Vn80NdoEPTIVrzj6ZhMtHiKn3GMZqHJO1P4/t4i5+TyCLpt3w0qii
LqOey6Dr9wHdGPb2OuTHqP7qt0Q10PR88+0XaUxyD6XaknISB/gQZ9ZYZu1R7PWAEevW+UAvys1j
Hb5zPkxi855v9Slk+jy8C81S0PTE5RTdOC6L0sDZtDw3+2f5PhGWiqVwURYAvRlB6/uV6Lx9vmpH
zgjDUvsMY31ui24mLkLXVMRRk+LYbhXiIDJqlylqI8LWaYVKOISd6x3LId7Wyy8iHvQ2SW7/B9nd
O0cKU5TJeLCAe3Tt7mhwqIJ378CX0QJL3UaHoyVibEGU0fP5EiiVC0t1w+zqIQtQV+G1omFxANea
80jJ7q+ZnvStlJqCwePMgvl56R1+S+1sDip7swe7VsEiFlCpsGBpjtWluXGNiSD3ZZEs0ibSWZeU
zlv9Dr2fJ6RCVVfL7Kf32mzSekRuTnzvbCfbV8RGGtIQVhsRxQm7fgiQKKbFA7015V+q1E1Vd2mf
Dm6AfsEtXz/Es0zd2JWng6vk5II1wes4/F7xCdG/PCSEfrk1fwydkwXn8yUwX6SITWPsZiyjjrPO
aEtzZjR4Id04gcz2LhbY/7UAhORICgjx0GSDcC9NTainIh4iLgokjndf2gaTDN6YF/gPwy4w6qUm
Vx+1CiF717uImywloFZSYXdruKPdVkrg8HgE/pzhTORunKN+h3tQdr6Xqi9aKFchnDVVzB3QIinw
ReUBE0lNJ/bYTOz1RpDs9QjbNOmAaMePC6z3+TRBojPa2po7N/Ajldu94m3KJ6gw3plCjgMHjNtN
bDiCryv+zBMO7yrgE7SodANWBrGBvK8cFSBNkJWrl148/P4ToKh34sF0KZXbsNbTsJ+C4VLqpbuz
GAhrqeN3DOIJ9cVj6ejBUZp4LBLBRTdG463qm26NoO4MaqyydYjG53DPeqOyAzzvSfRbapA1neUL
WTolvkckiRRFfBo/UluEhCqEYYzmKb/KDw+39y5w3OTk/0d56HksXLEGD7oL4aTWKuU3pdeFPJ6v
Ffia3mxFqvQUxa1v1pjm54oljKsSrhkNOii48fjV8n5FF7b0pKATFcj1ujJ98rfxXA2tmNWlMKQC
NhRy3TWtRlIgGZbJE3zJ4gZ4nxn+o/meLdUd0NNWN0zwM4epvW2pwMDsc9aCQnQMIsT+begBzK4q
e1F3t1dLHhxs2Ew9PnP6t7d89Uuum+zKddg3+HbeEm/zqg4Et8dDaZQ83Y2kb11LX7m4PxQwjQ9D
86A0gb8VgbDd8dJmjKE7ZIdu+VRsYexmOXaGpgJuvqCByz7yDUlzR4Gbsn0ax4dX94r4Z6U3NVFn
ULVXNINcwWC+pQr0b2TH5tWU4aVeR4k/fEr3hInR+kSuie7NfSK1YyLfrU3c80gAcZ9yCDnmkbCP
GAFuVXTjCCgiZ4mpAAzWHDJH0V7L7Kot6RQtX8h1lNLvUGsFVupwrB7ualhGM9YR1D48HRpV7wlW
QZCqsEwUUJMWvgKx7rEpzilWxGG5hzzGNlrtsr5bchp34K+onsNhH0OWffkyLMWH5arqRuO2Hc2D
uru8w7g7SO7ghB5cMyb6mT2Rl8wKyN+/Bs5xFBJjhlZvF3yykiJQ9cIc9/AKe7dlmJV4DoUiW9I6
TyBANuLnDs8f1J82WPb1XLce8b8zti1CzZwuGX5va2GmGBdr/SbSVRgG5fjVbtM7nrBPjOxfs6Zo
1+hqBIlLi7IHnBpxZpZx6c89AFL+ik2w1U6VYwEqDt9iLjW8IsLCJZBhsFS4pXH4tj0jE354sAsh
X5RF8jS5QxYIMNWw7f0WN3xv2ygi3sx62ilR5bqA/1uT6vQU5hqSJrwIFLtaterBDh7ROiM8KkSl
hO/WGRGNmLbN+Ve77MouBzr7YNgpFPHAVAs0bnueL4shJstfzKI5TFmHtnzblfe1ceXJwCrJFH52
ZErTNKIKopKWX/KuE+5S80Kq5jr+rdxCfCjtLczLh/23pv/r8DbxMmEQ7GICA7Fhyf9gpIPlC1Uo
gB4kfDFLdGgKZSxK/Qr3IuTd+6vyZyx17YyHfiB0Qh4hHMesKllrSbMu79slUkQHUFHFwUxu/aTF
iIKnGKS0tafgFoElNRn4zo0Bo8j4hvGXD4EcaZGlH/6LGhVzzuKl6kvva+zcQsAdgXiRyxnXIDTp
7Mg1GyZ0Y9255oyL6RI48HUymjRpXAI1BiGkub0HRIUMTZPqZL7yNQmWO66l+AmDiDlI97o917fW
I4OYUkylFDKmvHjdApQsp2ZszSSzzA5vISY06o6iODRVOMjMXIpCwknACiyyw2S6Wvbmg/DtKQBY
NTzLvaklmo3OltpLY9czQd8xkYP06kyht9ew+rj/epaCIm42AftL+DgPhOXOyo0+OqSFA/zotEzZ
6fkHteg/8fQRb5MysTxwDWi9Kou/DmoSb6Zb6Lnybys4qPximkD5o744dupkECiOO86hJp4Suzpz
c9c050cI+b2wZBvyFTlt5hnSapr+hd15iz0N6qbCK5PEoT5c9ueVsXF3z2yYbIxkgaMyiDYuuo0f
TZ/LU07kXQU5gxFWhdLFk2IzsLrSrwCNlzMYCCIAtY/qqwp1MfdK/DAsrxeNrDiChZmSXtUgkc2J
WtGzpMlPZ/xtC1tPNubH0s3opxBRKGS9QiY2Z8oLbQe0JEPTT/MUQBInPg+ZW1YfeywTYpuiqLOD
/j+uE3YlWTHrRfyFOrffKo2XTiPzsYadkWX/9FjCf97/L3DWZDb0qpQX5xG9DU4JdtB657V5xCDg
jFIXadovxJhvg326bxDdKD8eVg9a5wEBQIsANyNyZCBEjBA00vnWCFSxqKiTi7Vc2LVLDt+H8M3G
uaThexX2cTP5PsL9X0BJ1bPcTwsTUiHkNc6p+0hNXcziMj+DY+Stcxmz0mDYhe8ICHt0IS0g2k0U
nMsUoT7UaE53rdFQa6DgFGQKyh11eSX46HkzyRBv8fW1wZA5AfUKYj9akjaaNayAtWng+VKHlw4u
HYhZ0G58ayqTgdOiWnXe3dib3GLz1UI6cU1ogCODGbSl9y3xM1NunYwzxzgRwDVDyNsDEu9NFaAx
b0966Bi/n6XyMs0J3iqouC8URRKqC0x07BvqpzCUGHoGsasuB5F5lfYs10Q0Fo8yLyyf4YSKb/eK
72A8yb7SgjBy3v+c/2JwbdkeW5O6QD1CLlE2FzJu01+MhE2cjkhAf4nSpwAUxoX/sFZevEsXhI3t
VnXE3cTci1JoKLk1b1/QynOZ9CFZ0nGVbO28RhQQDoUv+NNeOICtHRI+I4U2z1rMG5aqdPCJjT3/
0sp4IXbQdPLa3AvvcO/+CBK9GImInwkqFpbFdw/e7LGw7GgW6BrXYIfJBpRJoFEfdQdfRm0cgO6r
9R5h6FGbia6IR3UDm8vfgTViGzAse8ZH6Mq9Ifc24wHoS9VJAXufr8YfX7q59dZgBP0m22Ibg9yq
2fwmsiTzxhYHeQMzlhA9GpEtmWE8nWV3elIqT+o85aAkoh4uLAssba8aMe9EmR2V1xAPAhBroklu
U4oqqFFWZbhhYHCmSVr+/lsrh9IpUldOOdC64imVZBw96XRfWDfbK8ucTSYMWwWFx6g/DHA/tP31
OjIhgY6RDCjhmTOxH4SBkI4LtieLsnj9iiSrHgzO85jjrzuTMlQMfrc9uJDjf1aKOBgYUmGyRdMP
e4MbngW4HQuxEfPNL3wVC0kOqy7qyAxoB+YjHRIGgFtXqMt+yLQXA9M8hJci3g95ZDaoKLTXfE2p
F3/+AEvVcZDKQwddcvhF79z/l/OQkdtyXL5FCuz7Hv5F9QK4aypH4cFhDq0h0F+ryTE45uH1VJx/
P/LclBilbcd2IBzCJ4WClofOXiuqY5UCFCQNTUI92OpIp4deElzS/N0zMUN5gyNIRvO8cf4acO3Q
Xjnfr+FN+1xloPQD3tNKJwtYSZTBG4NUiiF9eBj72h0lIqKl8Jep9yA3j/ectvrf+Xo/T9reMEB8
Bn3Bn1dwpBrn6efq/Y4FdvNWVfLqMOK7BBWxhOcNV4WtlQB3rVAYCP+pKMct0tVIO4o3ZQtQUyVk
7hLf5Z4SHzLTu5Cud0RIMu/MuqDlIZf8lgBUUss3+QAEzo6b2nXpmTNNrqcZb5JkPZZIEL8s+N5R
09xV3V3q36paLrGJw74wGocklRu1tdSuOeMfIwHqFJ9xkxAVerYP21VSucXqYuTQJIwFrQ5nvqd+
CCgyoBfoF7xc9Njv7I5XyjbQUfJ2aX7trMaNwp0QLdVV0dpVTE8q3xvBVIiBt7e76ezNWt4rXWaG
T71SeW4Q1c83VnuwLUa0zGeFTsH7MTk2kafo3+5wyMKDjq8za5rC8+j9qtuRdc1eAAFYshvHPZwz
ZJmD3b2LJIiq79owCqNOiHn65N7d2vR0JnVlAJSmPtDvT4VH5A05WxBDr6yFmQstBbYixwXRAq4k
5p1wu/161Z5RYCWLrK6utK8VoOK8oimq/2X6XhYltk7/AhKfd+3gAKo7j0fAq1iliNyUffpAfaR8
Wx+u4orS852TgNMJGyjTDUYMa/+EbQfZ5eBZX2L+Gu/SNQ==
`pragma protect end_protected
