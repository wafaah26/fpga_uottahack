`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
IGNlD35Bzlvm3+YvWpSY8+LOhc7XAtL7YRa2OFGLxwfqFOoiajFV4FGpmwSaCSj9t6vaqUCugKqJ
4cSC4bxkeZjQL/mwevamzV6zq2cc378/zQ4pcLC4lBmKsZP0qwZPf8CpKbLZMPtxsonVhZS0Q3JH
mJPCg/PHiYBmtV47mRDINHvMOP4Vy2vYrR0dUZZ6A8/Bagfuslz4BQRY//Ii3VYeQo9ADoT+Aiir
mNUuoCZNhs/vWZj2yJtx/rq1qOfySK2buPkVK/Gc9MsnOvWsGYJHjChjiBVHDhjNPhisXMk5f5W5
JoatkqajjU+4WXlHCAc2IljCN+agQ/kcJrp7BA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="Z2BFoYaUs1+nd2RrFPYY3aINpw7vSpy7vS6DndfwJIo="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4032)
`pragma protect data_block
4Nb622kKXg4Pd5GP+nwMv3lLbRTxOvUhfd++hVWqqCzOpBwLMg8IxwYiIqR1z5DyxP0QHmZ24kWv
NHc1TKgejTz5WXrw9P2m2zaH9uLi7Wb0mxBNjhaIQ1mhCFFCkWVxAUYyAm+hI4xUAs1WWuineVKD
tym68Xb8+VwfhFssQQaNc7LrUcfNrmVTgR8LE+wGvcgJIPXYbVtXz4yRZFN6ZXnDC6Y3V767xbWu
3giZHiUhZaM0G4DWhNUEdqL9U+qVBJ4WcJOijrV7ZRxMomOAqBijJIsqq0hkwbEu7977JMs/5ef+
Qk5x8GfOxf8Gi9AnZd54iHTLvus2jorChffa2aVBduFDjov5u2FMOQDOf+y/mJdUiK/XcvqYt/bE
KL0352kK/IGuTjPs2FinA94cfP/NNojYKUWLPJhZuo4mMOfIMyr6TjTtMgXUvS3eFLsh6q1lRz5n
WTC+YdQ99LP9n+FcvmG1I+UV4IPnGGY8HX9VIVB/tqLN37mHWk6iPjUMxK6wpgpxGXfizMjHy4vA
VL+Zy/2jcHkqD+mW3RK8PtG9NLS38VXSQjdToPSmgZVtRFuvwrIscbrFkHMQLkWgJ+lFDMm1Xuda
5mWVm2WgNZ3KeDiIXFl2C6JzAY0mVMLSoPJ9RO7nZb2EtfGYEjHqg2mGbBO78mtJGQXlVURIdYGl
BvjRAXj6KpaxfWbEJ5AMdKyk81LZzxv8ZB3SastajGAaP5p7NYX+MHxkw3kumZfap5SLMhLQimGz
IglLTiQZF3lRLR4P48JiViLDPRQHQw8hDzkqhgKFwIqdI5o50vZoEp5G9tB+EQQV78Lqx2W+23bR
A7RHUj6a9Hi8EZ+wLfQOBuV0CIj+STZbjvzGjQn8pvvfnNzVUimeCq4zAeoNK5R0bdZ55+MV5yDJ
f0mOxQzPUxbHrypT/NHLbXy1xklCTMxKFgZtsEmF/PskW/U5V1WWCK4C6DaVwi444pxfBmvJK3CC
ikS82IDA1S4zU0VP3RuMzsTk2B27lb6zHo/dRFL/bwlrUIhUb/NpM8RrPDpZZO671mfk8r6Xb4sj
uRPosNtdfZsgYvMZw2LievuQknh//XKQSnXB87nNLgvnNf1Ac93mczJalfVOY4AyMqmeSZPX3v5g
7ztptCKSFnWsHNHkntHk24WuA8XMLMNpe4vZVFUC/kSNaPb2d+V8S3gozv5ayoswmj0FlA3g+Y3y
iXEZ51RKe6U1RFoZlKpCxMXqQU0BGZo75AXayFuraWR4RgxzXkPlWzvzVXXoCIf4p2xhAxth4B5M
Wg+uEbgs1SKOMwuZCT4YPuvM1G3GWQX0F8reNmgooQGoRWyIPrgKTeULTxLFBd30RPG6feojgzCG
cRRmZZ3HYYfpi+/mqFHbMAJ2XijqiFnogXWu+0X6F1UXg1zeiaAl/hcFYZv6izYPCpNQSxo+oDUd
5J81rR0fMV8kfeOFIPVRMkxac3MAHhguWgjijmAk7DwG8vr/+5QH4A/wWq+jxRPZKkTGA8S6Dxeo
36byyKIh5kldRSNtX/1VZJt0C6v47kU+mt/EwcYTLbD0sGmsxlWv7Z/0+0hkwfKZE0oz9a9/08Wg
bWRfJlAqmyGFmnHIKdkM8YtqTKxh3gvnYEMFDZYNU4U5D57BXpXlRoIBeYS1WEIkYT59FqQp3vyP
VnZxu/oEVk6O7cHYTFV66DYqQXCGNoeUavfREpG4P3VqPlX+DYrCeyBkcpVwy93mJsysIpCaqNm4
hRHfq/aKoeJf1m6iwx6JXbS2qlRZYIuE1f+TMlj36jbfVRUeBVEgdjW3L9A3bU4ugu43sEA7lPGF
gjanN1EPgxzkfG1MAvgLP4VDGnkSsnL/v4CI56mmLo+3yqCzXodWNC4ciz4971hQ/XTogbqprDz0
rkhgOqoUCGN6jkRaeeANZNF4tlWv9u668Ry1QVjo8bgbMQ5nRW61KwMP6GV9LXxKuRhOVc5KDATZ
dqggS8jIClxTsG4hZLBOGilbOGWvkhnLJSzl59TsAevC+pS6EA0zB5OXC4xDIRyCYs1wERpEupNE
18ocBsdSUzbDBwXABKW+CH4HL9Jkw3VduPUDRSPy6yUY6/IDmghyojUV8bUSHNU0EgJP2xOm/4bE
4y2FmmcQEpgUidgPrKE8uhlXCrSUZcy4PkWUVUu4/uVSgzyW0Ry56koCrB5fpemrODJrtp2XF3VO
YhWZm0UPNDu0wTsObr4n24iz4ybRndZKALWHb7v33fcX81GwFC9ndlqKXONO5UutB3Ea1tkBXA/e
tzbiF6KeeP9OYIs+aaYyyibnCBv+55/1P5nW1d17VzXOe44ng8y33ONU3ppoMQsMOBi3eU1PEFIn
U445yHeH7k4J/tpbO1GvqrgsClhRBYHnMDbhEfLJDpb0a4qDZM42TnrIViK1OCZ0vdm38/nTkdh+
HZM22j5JVXagPiXJenU6K78gW/x256THIzEJQEjI7T2OfRqeJNhpXQflz7QMgJkOTeCVKPptXGrJ
ShYKGKSOCEW+F7P6mLMdbvBToX/87fqD+F7gJvBMkRvDNDYKxeeVRddERdehpFq7GoUKSI1tNOja
PndlJo33acquHEkVaYuVyDvvcM1skgnIxmbjBRlDEMC5lSdILsQFqQ6VMS0N34rpoYQKb8U4nUzW
rECYURM2W3R2qexYkgOSxqYNrgt4F4wejQ5hzS5KR1eexcG3MTTDKJiju8Km1P4VZop8ltZTDrhR
sKGud64nG0SBGU+kVs+0LCiDTvklgTWV0QPqMe9k831xz1I1B4GKPSzZFLY/6AXrb0HyOGRlkrYH
TnUg+TI9WW8+JO+FPoyRQHsVVTjR260/be5KixeBQHPTeTjo5OU3LZWM40Jip8jlupEepWSCyckw
wNYJAZ8WZBb/TWexAe7dBfkhDJ/OppSE4BVhBWAa9acvVb1hL14XtX2gOALZxG/O3LVeYohCFQRA
CpYoW68Bo65pB012krefUg+Q4LazRFWWZ6TK5TjUeHPrgvJmeNLCTme6bQklunjfD8b5R+YMpN1L
TraQZaycJ5HLoCRmnwN/CbqIUWzjHlLv/nMH4xYLvxSd1bdow5rzoKZGTEHdOuAcuhJHg4LaYmBv
xt5PQEyLbXm71cz3RBo2bp4UmqoywRQK4Fe8YLXOSG0xDaUnlwun+9+Dof+gBJNcaB0m+k3ae8oB
PhAZtW/0gOFtQk/diqLXZUpK3ocu6eVzm6GjoFPEilM1Mtp6E5WorGloXvMFupZANi53hHVPc/iF
6mUlXobbH+53i0c4DVBcXvZaBoINdtz+tQu4eow6GNIbjwq/q5JkOYalt6SMV1SFWKBYMzNBzlOR
CHcZZfw4X9t3TeSKeR7fpXORcmDbWWCN8GgH2nMIDuMJOlcauQRxC6oUYL72WIbkNPEPAx58DVXi
43L7aHvxZi4xS2ZnZnOF1L5HKdDCnDilTCosjPkkgZFDIi/SNioLMKgycS6Xg0oa4q+0SAhnu4H6
d7QQ8xJXFLSrWerdjA1aiCyHSAtcYKDrvl4nlnsxJ+hpm6xypqiAWkj2+h40BUSccCtCtxHmOZWV
kvrFhQsez6ni2hU5K/778HA+MeRWjM+mqKswa5h35T41ozlwm5lw5QqM38LmvrPUQ0OsgqhYXtLy
dWqNf/A3lFHRKxlH/4bFAJwh/3YpTQNJPIU3LcdkoeO9Oj13rFbBFE3wUq561ehAdSTBk3CvvWUr
jxGEj19gtCgU7ixw8/eFquVhRZwn8Ix8Vha4KJtZN0uT56qz4cFgCP1NEHhdwQZTDzJyvCqq/xT6
ypg+zhHc8+j3wawdPHujD0cfoVNz/WOVYv+lJaLeRYs/X3/EGuEC0J4tP99M9nmJ6I3fB8qIZ8Vd
CqadoLvOfFyMZkUqxYOkteZ+WqlCxzyO6qLAL3RUlK874hV1pyqm6DfpXI+Ltlvo2yothqtUwUaH
60ai0rbM1EtiztKuIlR8oohdkRFguvxDuw98zfXjfuqlfhZn/MfZd/pYECNC696bqBBt2pJY0pH0
fpnOzN8d5eAOeMLcAKmWjdzRqO4VWpOgttkjhYE+vp5rYkzTVaOnsYhFv4tN62XCmESviRle+39f
6Eo14ElhcYpqLH9kVqFUadb/pmE9gw519EUB+0A+KK/xK4x9OQgzDBjWt+1oOgrWMqCuU/DPlbpk
WyLhM4kTZAScZwtnCboR7G3zp7SwI6PE0VofmRoXpx2why8ylQUwR31zVvc+SFt1GuuXBrodiQ2M
8nWHzOI7ykHGEUcBfnJyspwd4vyAwqYEJyTEABQV1V82URRS4lQ9NP+1XkAJSANpfTbNHZ/zhCUG
GetV02kwh9MuyN2Ykj6w5TUBbsV1CbErW1lsoX4exIonZfuowxN8rj725/jRThm1e55aFKr0tKzX
UsoItAM53e4ywz9abFte36qXI0KYdMVuu0ibQSx2vG2frx6NAGB2KTeVUqnKMXrlmtnaJSeEjwm7
RiMSvktAnNLwektJqIXsyq2jugS3muHOy4Ad8i9Lo8RuvRR+IMhh8Gv9L7ENA29cFUIDRSFxDnMD
YgClA9z5dY03l6SJqsJS+lSt0/Fs510v4YIYPR3T48I4i0vEY/XTmq1rKSfPgh3wK4CC1U/LtaCl
MR4U7D5iiHiNtqXQ2QzOhpLWfwvp+ZnU/Aqe3oOEMs6iztzU5wAQ72jo3Wv3IqvtFvFJr0c4DC2k
MAOtP3CDFk/46Y95b/+spJlg5pKL0amnPuirIgf6X6Jv6xS6i2zg4YiHEK2mLrzjXX26Zhg/4Xey
8y4l0RkZO/4Qtf+LIUnLnzQ6lzsK1esg4q5Q2Sozr+3q6nNXZ7vatMZYQ8rPbDKxCuYg/Npb7D7O
8s70lQMVkCX1ig5YjJ0XWzxrCsJjQWRxRCqMusrKCJIhl9DO1YaLEO1wvH1SAZQS1O3ZbKl36Q3R
8Bf2MEWp/f5pAOmAQchX+xM30y/j6Xwk418U20WcYQjbsxmKAZp60rqdneJScpVzw0uUZYe2RPCp
mYIy7o2905qTFgREJDKrFfM8nX4c6ZO1hm98vyghtquzYpy6swG6N4m4Rq3cwGSu2uxhp4tTapgH
TKCZABzsSeF/MvPlA0HZIQxe1pP/0AsaWQ7opkwTl4YV4nndL4KiGG4D3CMejm9i6Cac2+EVzvAz
gTHNNrNgWZXceNyoiCUPmtt7VlQDiBqr8MFLvPRyKzPbMIP6K/fdTA4rFVH4NVOiTZGOiUBjfQ3d
Sk89RqvuD1Kugu/gr/HIONRwNUMz32x9AOjHtFex3nXThyCP7EHgWr1hCCgWD4oHILvlv/JQjgy7
/l5ls9kSYPEM553Xh2zB93tUCu/D/yQEJmahg9odAPhGWtKmnHIatx2u
`pragma protect end_protected
