`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
BIn7YednpPAhJ86cugaRx1uKTeJY3SuqMIH/6pO/Gb+TNaVu4nRUASPOII3iR9ci/cpVcKZfQnqe
VvZFSczNz2V2Rxvw7RI7Jikf2iEN6sYaGymj2EaDfEFwhb5OD/CTAc5uyCrvOUNZD44e/pp1pSbo
/sfdNBAwZvFFFp0Tu+odkwW1QS2m9qGF22OQQMrSAy72JUAXzUNOOjpItr3J6mSvziUi9C7iSzge
O3gyud6tImv3C/v74pY09Rvc0DCqYeTxPaBKW/QcPfOmZiIhJeJoFuJm/7J6MD0bnN1hQgez9koK
y1X8LYJnHuC7kmqhg1zSrykzmVzOs4GkoIzt9w==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="9kOuRrnKbWQnIDMuYIxxDgqh8fzAKX4vPp15sCG9mO4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4288)
`pragma protect data_block
YFYF/TlBtIzTBCUwn0yxvREd7b2PVkU08P1EGIwuu25JibXuzK0ceYaKt4bUCclN6FQPtPA9Pis7
QXH0vQaBwOq2AgvpkWv5toP3Ng2ptTEYeld9VSRRKfEqauqvdSBjZLmc/c2yzb/kmOS8UOneINWP
fHS8NOHBZtb+4bWufdtUEMOFq+uGhqFg4fHZ7NZfCzwWbpXeDxiapEpnCJhbEsCCJRZe2frC+I+h
zQcofteh1eZq1hGMXENU8zLvQWoCVJOC4SkhdwpODpgQQKcTtRN+bDas2MiEAytO0JfzOYsLTo7E
0n1FrS5G2+E02KIPprTzVXO19UmQtzjQfhVxiGbeK8s5nT1kou9hU9tEnZB8gEWtSc2QefFzKWCb
JS04/j9QXbczu58BIcaOAfjd2ZBYLDMt+V9fOziWpE4ZmuhYrt+eaX9nIcloIDPL7BJhVpascmKJ
t9SdMRbXA7zikQUKbB0Zp9C4+nIlVuODffXvILtI9p6iLaYJbzG4EO5GAzEWYvoJBt2eb3p+1qru
h5F8CKGktTSSs2BN8CftprevEvaHGhv/0znjndN8SrgEF9ltvtX2ZreazSf8/HeBxkRGjn3ldKNv
Mt7gvTXpsX90gdLyj8CN4Kj1b6Wbn6CjvpbP1VOTT9Q+90RxGAvZgdwvUR9E7U3j67IeEAkZEhI2
IvW2b7tbwj7u3H+VWLQc6WsyxAHRUM7hh9Z2aJHLJg1R5SXJFIcl/HmaJGtHn8m+GO7aMI2p6PeX
LOioFq+1NZxGYhMNsDgGwS7NIcC+yMnXI1vEfvmMFGgNLL9GAJs++y8Xjh1EivFJCKoLDO6CLer2
S4b+6UQK8mT4oPCTOoi6LL3A6cTO2YRmdmS3vUsR/AxZ6eRxU1DgrCiFIuYoRawZfidfg300ebYA
XZsZwPMr65uS5ZVrjxos+g/Sm4+5fgx7OKjd1wbCa91HEVEoiS9pZ8KsdcnoIA01+oW/PybG1HuZ
ifgSEcLv5sTf8pB3nH2KjQpJt5CquIbPStWOISifUsb8T5oL7I9kYiBx/jzMt3FeYfyxC0i0mfTC
lad5W7YCgA7CTBVvAJ2tj0o1f0SzvLGE3fxFVFDnzOmXHwWjNkiXbKY0VaZsZfNBQaE/rg5/mhPB
oArAt0olQDpRT0N4SX5ollSv4C/ppcjvytrm/S+LyXfHa0Vn5q5nDdvnPYlvP/8CFGlQxoChdAh5
3OVL7F34jSyx4+Jdz9dCeeP7yPCqssn6yh5crIACCIFVnkkA2SbDoITo602uXrtLmgi7SRee0Z60
UpG3QbjGfDW4JHnwHCBL85oA1RzPWOq0k/cQ7+v9jSgljnekhV1UVp75ZNLkKspFANV1SkQn5MJL
MrCS0rNkvRywnSLJQzfSKiEt9hgPUiTuhYsSgiW+PGhBayX88hqqXjv/e7VMp2z0Fy7e2BrID2Ji
3JfVkqHPzkarH7ETE9U4UmzuXF/LXfVbKkpKpkHsx+7IMuayD6VDMziT5e6Ue+0sSLsUyFzXFKmP
jpPxd6S2bkRQsbPMefdaV4eNW/YLoIc+QM7Rx5RCPhp1OCB5yWsEENmHxsBNWPtqH3hWjH0IoBVU
gQqCwRV8i5qtLYu2Ild01gBDQgAca9T9/PDmmDN5LmrWahseMnm3agzYwg2IzaD3bUxw80YDoOII
55B9+Ntkkthl0AjSW2iJaFP7vDMU2d8Qli+XoWcGMsMsJGRyOuYU1DMwQf5/xqxoWwlRQ9a7Nrhx
0NC0Ve/rCFYrhbe/Gw6eIckFxiKz34lfnKvc8MiXraBnUL23Oy7++X/bHlrpFEpfXfm4VnHpS8xs
BOg0akvy3YqZRohR9tY/QX63wLlIfKIDpBfVqt4yGlAuahRSjx32HS/3kZi+8dXIdlas1wNiLPZH
LrU+61HYWr9vJBOF54rCzWfIDXVONY7sr+5W23btYzwFgllLOxsfwGb/oZBfljZGY/dKEt9mFtrU
6CIcfq3P5lLqBZudekBlnOOaTNcULNwosC4QihHeL6Sfx5S3HMIWuzuz1DGFfzOxnDjXC7AEKzmJ
83bQqgVWpLiLmiqxtZ3y2aw2rXR7X9CsijN+2iBNf5mtZHigVc9Uocd1qWP+79WqRKzxcg4KP1vn
Yt1XAepqNO+H+an4KYPJzlhEfjJ7OUFWEnJR8+CK5vNwOiINRhuq7+6Qlb0jN7VaiY54CVnSQzt/
/GKMDJOhS9BRX2pJnBd3cFQWzww+SzapBTNQLo8MZxFIDLY1KhmitUr5SrPQI8XRxCIc3rtlZQtm
FO8BQ4jEO4VAA9et4qV2cZaAh7sWNqC9s6vACDmWxJJ0sY22ZqislCNRwSKyZBtMuZ5NZHm1EDHE
YyoOfw+9xppbCFw0em1wJdTmJLwa5PsOFAO4WLwvGxU/HV6ugBeRQUw9Oj4XFT384Pht8josWc7V
+gf3n8y23hVB2oN5BdHxmOWSJDuGmhBheHnDsG6IorI09KxlxQ6XkItSYJKa85n3oGZ2aCB6D8iq
ing+KrhgeDKPk8WST5+OqXW09k8gsFlK1XDH9veC8+53Zt9RLA3DkRN2CTRCv4618YdEBEJxHL7L
qg5gTx2ZQRM+yp/eKRO5VDKKCjKTVvGZd5/VMF4ycoTVNiUwXTbX/EKfLcsgbuKh2oQBXO4EPo63
cH6OtuhJzJ66xJ4AiE/zWZgLYbIlA1PDEd/UtU51L95bwXQy32I75xS102i+cONBrunAdyu+USt4
uVCUTL++vSkKGh+H4KJlyzjANvb/hxYMnL+4t4bahdgz0ntwGmZ1Mc3aAlnKuR0DfQFtk/HnnJpz
Rg1//7reTEHi+aMYlWCGAD1rrX36CIdJDNh8XSfptqM3j0uZtElwuyadYDaJPaPxvElJYxfHg5/A
45OPDdWsNHx9Q9BqrHQh+KT/OiWmmzOua60e5jU1gpdGaJZDWaFA6rTDifjB9ceVBP/8B+kUWG0X
Uh/zmM8nFqkcB4C/4OaTwHBycrDN9ETTGFP7+w1hro441DLyvyiWfdTsxFF7sug1lUQc862YcmGs
uLbkyu27xaUmdgof/TCnlrTohB1JPNNpgMAi/kGK5PcHJa8sHDp8OuzqffNt7Zi3gcyrGEP4HoSz
ViNIsaPRLd45iAmjTlmkKuBV5xsxjy/02nB9fWVLxpyWhyOPwLkNqnJeU1SXRZeNfUok2zPRht6X
au6FIX8poNW/BTpdj7Anwp3OYu72dbpdB4SwMGWi9exXFX7YgPZVhf6R19xL3/IqDIFpVN+la6xk
BhLji/lgrlo4rxtLTLBwImBmOPBSIxeGV/FcYWUF2aZ51WVvvqKzBVIOVcgBbrlWk3ZNqad1pyKm
pOTii/tih4iULx1PER8lNAEeL8Z7703HQwjg709gt3Z+9S/HtTxDwc6P6pzoyrMP9q1SSumigOHQ
MBycpKiqYqTr3nF+dSr1/L4cPj6gDYLeOXiDiUQU5mWgL5d7iwy53/g/mpi5zBckhRziYwOqi+bT
O8VRrckbzUETf3JiTHbokwLc6hPFhsShZQ3T8Rw9tCk+pqb5XWvanSdVDyM9Tats1UrYV3chmdn5
JEGiPFoeiX/UBe/SCd+Wl/csXxsUzfQrC11e6zHGCUwHcDsTbgDO3ZVSYalGzGlPSPTy4SQUkt7w
D0Yy/Sr7S7yWH/iJ2gKwupj4m7cAnZv8GdFeJpS4ptjdyjawEn34tghoqTeWKccq/Af9sDkww1HD
WTT79B0R16+9AbN2jqJbPAp8RP6zKqJXP4iZT1Yb6I5EWNTDWARdGvwsmV3oPtUmDlEAsbSE5XIL
onWKS0VcMaFbX0w5GXFYWA06I0jGgorU7KMWgvOjLPNT/juy2CZurK4QBhy7WSoQe2KIBTXomjph
zXXh6pz7a0NkJHRmOdwajbdH2VCO/ooKnWvetmP8N8rLEXL1CPjliB/rtgo6OBpO+HT0XFo+99Hc
C8jAcCZl07obtx/ei45V6s3N7iBHf1/zBfP+Wl2w1TubEZfHdTMi/7pjsar9ae9JU1OoyKVZCfnN
ZQ9MDSHWQJ60zCluk11m6YzfDU4KIVTj8Ja5Iufpb8WdCN8DwApwi3nIloiK+1PShcsNkeYWrOQt
Su9nyqN5bKYRL8MIn+TRqFxm1qbTj9lESublpvJsSVDC0JIjzVh8EjAEywnuOPDXq+dXWWlSCwZZ
uOrtAhpUaLEXEs5rUkN4nM5BZBaEBq7wKHWeKgD2o4gTsKW+AW3axZ0oi9F26pm8ThWSAXtDhlt/
hwVIOSrC42EZ/8rkbJppsAtTTmZn+6u9XRNmWoK3Cn1gQy6bh4ENrXumv68ITy6sJEcHWJ1/WBv7
og8eTR3WKbUMprLrAiyFyMjCvvw43uhJSzDSKSzWsHv06YZ36w2ZZAOTfmNB1C1jM+lSLjiRl5vd
AneiesrKCxmFBuE1nFi83NC2PmHFKQk3bWE/AMrWMl9kC0WmZOjej6Sc1TDrNNCRcUUZ8RKj6IJ2
6gcR05XMJ+W6q9T6P3qSoX6hYxuEfd/ETnqQocUfyRvuBVETOzwdEfs4RtV7uR1azllMyCyQHK35
o1vHCTZR24YuR8k52gOa8a6Z+La1O8JSPN1nWfF4byHSLtSTOHYooBc97sdY+yPYaBZ/lOvZRNFt
zaXtMWOhgPzKh9riyu7Jpcnf40YRZUkcJGui7w7psKfgGJRNxlTe5GrM0KEj3ume4ijRAPy3k1AF
7GXSDwh+xXMx0xtNyDIpy7J6E23AqIuSv9hQnWSjw07mvx3TPBj+mkMlWcPb34qSKxprd/VVzTgX
d6qJFtUPDmRNoWzwn2YjNqWf9E1PzQYL1rQeaOChR825Drbk3TvNDXiiF98V+DInPE/N5rj3whHr
XkluXiXceLd6uCxlYs1G1xHDRr9N7E7GFVQrMIjb/QnDgLFqSuYGqGkRccz7WHcr6BTking+A8j6
/IcbzkMVvdwKdK57DuE+827BvVnnLYrk8YeCm1ylFDF0Ueh9D1mF639ViB1nLJXwstUFgrkepmEE
QG8aScV51Bulayoj8U9cdmaFxdJJaAro09dKl03Q08ycxRH4jg8vjTd3D8ae223bm659i2aoE830
48Mxpf7GuL1tZHGZLBNiwN+EILTJvl9ZWlJu2MTNDDXbjKilZRupOK48rt6YR6C8FZtw3LegSA0n
9dFCqkF3IA+vIg/RUNJirph+pphNi6wylONmr+DFGfHlejXcK4AMcL4pPl+RbDgJ3Y5/d9W4qKga
DKmqm8QqNDwV3Fb6t+fjig2zXhYaa/wI64mNSL/tt88BOLT7hl68HnXLuIeiBodUBXIYx69d2aYJ
dQCrh86Mep4ByKB3ziloGQb75+uBbrb9NKCAhU44hCWoTrK6Iagva4W4yCo7QOQ8udxqeLcg7U0D
r2ourOZFAYZ9N7BUcirt2H42E9B21EXxbKvxXjs/l7snY6BCpSAHBR4SGN2tMUFPLEmVfgove4xM
XUgM4jCsZDiAaE0S+Se8FC2WY61fNYh4IE1KYM7EHvTQ+dxoiMI6G0MO5YIQe8BMVvnwYP8BlUQF
L17SFr+WLFqrTtn/lSmX13V4QtmoJpSFD/AuAPn7nmDwTxM7G0z0OJB60QG8EC9F9MdFDu3A6rdB
xnusyia5Hw9ImnB4mvhc5b4RZEqWZ6R0tE11ta1C6LqS9OPTkcMWWAWtlest/fKkE0c6H7rQaLPb
EM1QRjJpwWvH0xSp4w==
`pragma protect end_protected
