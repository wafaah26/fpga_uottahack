`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
Xe92pnLAzIYxdYvEyF/FsxxbZHNGDBjLzajE7Y3DBsB0LJE3o39jQz3R+W/P/rr9IE9VEiPNpJYO
ic1XXH3/emD+Twj5Jxce6+JNHzTS3iG2laJ0L9a29mOpehHP9DjnVJCQdIFdIbCXoqpMOC6Q90zC
M//CzGR1txYFfyHh4HDG5Gk08P546wPHWybomBsUugWH0aWux1adhn3oJu7VT+/lV+SFQCFheN5R
zFXmPLn9/GKpDp3Nqn38Gci79675/VeHMcI+lXIWQfhSGDWVyggkZxw8m6LUh63aoCHOen4fiC/c
YxroKhk1vUTjYvNnomYIKHEtDYU3i6w84tmVGw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="8/rVXWcKiCXShUcYJav/lji2RUduwoQYqT2UelY+4u0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3392)
`pragma protect data_block
TJ+/80viyF39X1pjLPeK52XFW20hqEh0OwoQty0H/s8Y651bBZlsBn/IXTvIJzDzUC56BmD6R0Ip
TWyS5Vv2iVBe0gvQH9QxXB9fUkFd4xL6gfVDiWUJUT9EWnbAY9W4pC7wla5weizYFLBINk2W20IF
CkBQxkSn8iAZ8j1p0IcFDvUADOhaHB4gZ0LllNScGur0x/5Nfyr5izpAsmJltbE+eTaRx25oK51r
BCNfU39kJvldVa0yYYl0DcZTji9lecp1kS7J9NWjBg2yA/MHEKjRIiK2XSUkRrv6zWcW7YrbTusr
gZa72ygF9w1f4nmViR3rHKHZ3H2HULoysHsUI8behfdCbf6SdL85J/WT6+ecntYlzGJ7VLfUFLxG
fS6mJx1MK3ODNv8Nsyeid08VtDjLmm6O/DMDVVN31RgEw1JXjeIb/V5krXvJMYOlvE2PaAwGzTwn
WmX2VugduwBXAp7OEhSZdjtAcfGfSe+acshcoLHynxv1srUaGLPwcqpb1b1chrsg/GGG25wjTm1F
jhuQvxKbL3d2V0agJlXvvmq7NxSNJxVDmV3jVFADPfgQqmWOG5Ip8JL4p3c2sGRIa3u3fZYYmMac
+Euj52NDjp9Ff9n65x/b3gNE+7i6e56GoqkANh6jPiK3/TZAlAmLmMLDP9jK4MEiNn3eVZINhR6U
07UvoacN94rnEbFzgGYo8QLqT/l+sshyermrWJw61N//ls1HhBOqMiz58ICF3197MdGkcjUz3oXS
O1YvzBnPCxpF6eRzGDE9tJL3Lq81Q5QCBj1GTLJNcW7zJLr8aUWEnPAEBhoK9Sx5M+W3EulihG6I
DSPqVVfFqo2vy6N0PwSMrzlP50QODGWlUY8w+JLD3+e+/79RvE3Rdc4LOxCedlh4mJay+TwoXDLC
I1oaIKxamGlKpkrODUkJFtVSeUMWLtHX8i/ooj8qNIOyjqf/bvbvdhaNU5fvkx8U6i+8xYuqc18o
UulOIgcBW8Mbw6a2douHf3R1iYHjSKym6twyDHzwLIG7YdMVyUXC2ANCP2DDGRIfbajlsUXs7mma
eceOrW+SgQ/qPCLaBeBp5xP1e/CcpeM2GKDd1XF/toUyQz0qb+X9LvvuBtvxQQPHsm+w/5Pb1J4J
uEan8pf+Wn9uFFlgkKoWa2LyDX4tsa94kN2KaBB4YTS3mroRwvFfcdYhZGcFoHj7eLP10ODejZf9
PdTObGYPupd7Ye0qIwCDE5CuBAcYCFDPzpxL7AGM9B964EvxBxr7mhjor1aUGn7v6k8l3ar5LZFY
OAloigD0GDF8jAwv4VOzOBbtOcBVR1L2F8itubEMCRLbCdXGBzkarM9F0yNJH1FN6U4K7vLISWA6
yYo84nM3qp3fbqiFVlxGN0t+MIU5/fusw/ruMNELB2CR8EPk3q06rpwIzjEMkc4hueYsz5/qsYfI
kY7zpdoisf3hDClus50q9J06TvYWiy/2bWr/cLFQg8yzDYb19vLcu8SGBuMJFZ3YjEVay+ZbVFsw
GpNUljdnTfhsWLdK9KW7OfK1aouwGG2kb/BMrwjlkV0CtcBjNUqAoWRR9nP0vr+veF14jeTkh0T6
F33ioxgci4L/a6Io9Lo8Ds1//A+YEIyh9wKhfbX9ZDIb3rCBjNDmJSUwGgfo9aFy3mJea+2AOQgW
KjJhpmAortzdsUqA64gqKjwVLvMdESJLyOttKjhw8cqY2DAWupDVCwhIQOvxhJRNMDMhifA2/PgY
l/ih3rX1pZruka943Xq6vQBSacwNiQE9EGg74rcmot/ujDOkR1fo6q5AytAXBY+kK3Npw+aYJgQ7
JTs02Gq9iDUCtqbH9dbd7GxO+R7RkOy7QX12GOeB1N6WR2q4KPc65Ws3acXjtI8yk2FGtfFR0r13
Jg87vBCP2QIAFBElZHAym7yMhJYHOiTV/Qu/4ghD7XvDKlyALN0arO5qQ2yheTZOORRM1Bw+h0Fs
qDHp/Wgwk+k1WBmJe+eyTDRpxSXM5B4iUuvSJ+1NH8NsvReCMcEXSG7bY4LOY8VJ3xmbC0VtPwlt
e1/TkD/Omtb/tZkV3ke9MG1kVmOu71aVXQHy//SUWsh9yUyJCaSIdcXWs4K1pFiTZ7Ij/lnZ2fmy
bpejVxqC7QsnDd8nAo3O1qNHUT2+1lwu9t6wijhwTsXYIdki/DTCooIaPIJ55dDqEDMaKA9dmcAL
aCdZVJusJxO8z/MxfpQH/oyZasXcukCwdfD29nYXYmsdp+MhGEk4xUUblyRWQ3LqyWPg0uSrSyZa
G53Oo7YSPaJ5kr4LuId3HlJeMB6HlvcFBpulTJAe0stsaJVxGhya0bX5Ygz8ZyHnIU8RCLa3sXcv
ofQeoCZuP0dATCX39psgHROturwIINlCMgynT1cGkRBfqNmr5q534RaxafgdbUDQhX019G4daRMf
nm8wrakrC3LIYUwEYgq8NVyul43rzZrlFUQglMPTg3/hD76dU6/mW/8mpNaWHwoel8i/JInyHnue
WPyUCg0Gw9LrDzZTVef+aCnHjuXm/uIoWjmAZyW8J7gX3IRpx9xzr1s4EImQ9Re6a6hh+Hr7dodB
FuT0RhNFgO628vbz+2QwSj7/HELgGOTaDvs9qhlydLx+pDpK1MeKVBQRS2FQyYingN/HkoAtOoHg
FUXcrHXMRB0pi8UwWS60+YErZhkP909zgxEsXM+DJkHcbItTqWIlKZRYdZnyYUr1axbEiZJFwM9u
sfwjbk6tGsU859+ltdTUl4B+wN3OnrY1Pm8tm14gSSq9yVCXbt6ddoVBh12JJ9+PhcIpCQAuua3N
PtseHP2V/27Nwr5CF56YwmR/x/ZgSda4Sema13EVhmK/K/HCQw+sp7kkf9+giS+CC5dehsNTRs01
w0TLUYMJwrRDl3h+9JNlDpk1M/byr/pjFJmrJyhzeb1lsTYJcLKgXwLOoXeR0Ta4gg33+XEWJxA6
vM4eRjalldDkGY7gpCnbczYnN0aJ5DO2yCWDuqFCb7O3ejmGS0VVKY1nMxIQTMddB8wHR2QNz/Xq
3EMhep0jTk3foOLoxUVkEJnVDhYcRpOhq+0qvLJn3G4XiiCR0gaOCeB1eAlmmYFDnSkWy3fO8z33
uIKqdOCDJZS4tVKd6YuNSIsel8yQzDrXcMHLFp9vim0HYQODW56Yg1VcdeCkyysHE7ybdqt+Jx69
+aCpNO3fuJLYaQWPQYNwR0EMT531lRFdV9ZQ8ekgqbrN3JVgNN4UCIkMLtGZKKhni3SBuwN+zRTB
XXzfOCsyDJNlgwvoZJh1W3oeTKI8mL6lGkBKLTMj29ZClXP9Fwz+TCBBTK3G8H/Y7I/G9qJpFa0B
f7IuvJ5w4Bi8AVAqsQkJ91OuIc/qGNvTZXC/wYZuxVj3XOXoGZJ+8aZf6DLuPgkbs/pKm7xwExE+
AY43/Yo1SnXbjmzj2QCVyUQTQXtxPoWHhGWhTSJK+RjBCT6yFyLdI2U7DMINjDnGAaZ0FlgIhu/r
u1NzaodCyxuI0b5aOVFJRpAfxPoeHzRMhXItERIbQ9KK2Oy49i5qomHQLoqPo03MOjjaECB//TD9
9HpQ76l5uvrTMK8eN3O5V9ydJzG0vI5zUBHA1bntgnia8em3GqJMh0EihlIZtFysUeX69AlL+8dz
bHCvs4uB/p8+xtf9VN6+Q0/sLcegJmh768Wn2CRHf7GnkPWprKReEo1kAvtI8TlKhcx9+JAUdfYw
K5T5ELben+BctxFhBKEiKhif88PP5dUX2wp2Rh1XJ5fN8raQPjCM1pqXAmVHzS0wRB0pRG6ig7NR
U4xmXBJJMPkbKV+y/Ik+512aTbXKafNK1B+vm7ZiK71Yai2XxdlnBjEgzwjoASRBUAYvJQqWu4JH
8nynu5aIL2bH1c2mfixCVszgG9SXeA7cAnsKCYA/ABRYhkA1sAyA4rP2xTbb47WegwRnC5cAWdrp
3/RMEkLGWEsYAZjgKE5D/QpudfeMvnfaoC0grieHatLGXbXvnmy1jlilggTeffElk9JdCokb4Krg
36X6fGmDeFtehLclB91+Fv7Ozpp9wXySVFNsBOibJGMcPHi8iWqimnuMJgzBbQep0auDhRGfqoVu
lDQfBdRarQh2A/FttIDuefrCzOSdFjKLGMG0f7ixHTcm4WT61AXnrMPjYU1j8v15DR5uXJ8CkEnm
nGAWwuPTxpF8UvENn67me+n1fuoPdV1TaLsm7wHAkh/kfpaDmQ9FKlYSF6DAkROr3epqQyIJuV41
PGfctilHN0pEZ/0HkB4xxdGUPbKe7bygKWFk/opV89N4VgWsdehHfhvcQGMzZx4wWyy5PMF8/fhW
1le/1x46KK7fImq7zfeGH8y7rwydaitqoRbPf/LwTkq1pEc+2aw9IKWq/H33owNxriQp6kXCftKJ
5sHEkKrl70uGat4n1UM3EpI062TIzKxZdr5xL7a3YCcWJp50E8afQ9HO+Z6cZgiPaB5Osl2gVrhx
H5V8BOP5hLTwEDxSeor5p7LiBRhb0ZOEloLNQsk=
`pragma protect end_protected
