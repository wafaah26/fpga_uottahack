`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
E773cKcP1uDDFspCxy4ynIbu9RJp8VmNhMQ2eBh0sD3viWmy/Hr4C5nGTqkIjLjGjmgppSV6bSYH
bT22c2IaPdRdPGTLjxApt+ephkQyo12JDyFMfgww5zd3200JykikfvCkPiowawz6h4MF71nas2zp
Zr3NZMXQ/4JkssKIwVb3E6dHFE6nmlRwXcu/JwoP6ggknZ5KwmFv3p8TNvZTDfOXkkZt5cFw7VOb
ig0YiNcFHgGtI0sONHNrW/IPsrECmzMal6461FdiYKq9qwjUNXCZ5zMufOmtuXBc1Hl+i5aZ3vi+
vyNTrwfxQFY5K9mICbTdjJkPqqIUmq4YOowO3Q==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="n4WNpMyj7AOqjvYCa1MlFnWUcDLol6IjtWy9iRRRkhU="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5136)
`pragma protect data_block
5loBdgx+9z1cbUPUgeb5mIT6qdCAqzmb7x2Ez8qM8yK9h+nrZlVcirqRvuJ8XCUT3vODeuAREMRk
tca8NihkeMdr806mr/LTcWhoJxNa2bRtOPhmCr3SXdWJtemY41mLg//1IT3VkrvsydC0/Ius34wt
aCrWIyu7TD+s9ad4uEFYqTD9GRuNTJ2QgVzqkmjc+CtjWSmjqClfhwvysaEB7ZQJRTzCeZpgOEmg
i+YM3tKPS8TqXkMMEccaZvwd6KTDgkJhCH94T05/E86FEQUElvwNHHU5Ca6baZdDzvqO4tDJW/9i
qBIyNEOVANTyuSduTrjosdP1AuqH1XF8Y2FEsM4WktvqdrHBYrGusBccUvE8OdKAC9h7qs5A0P5y
xaHfYTG8ykJRCm4FCbEBkDE485aOpC2TinclxjwDOmIrBUvwOrbD1QLqR/0i0qM0oTTlBUxYIE2n
fcsGneo/aSZ3mA8G35z+jrwYESEIh+6w4+MtthjaAsFCixfhtz+EYBvml0FlEeNztwghzF8GaELb
N73oU1I8JarLCZqMkSilDd1yhFJSL/Az9C80uljgHa9GHzFxtgantVRSaVAsMTfIgi4LWFSosHo0
YV6S1bYIaufQ8cgrB/Mlm40PxDE1/wUXnMCt+XER1QwnBA3btskEcj5KVAbxOqVMrLMaSCfffKs8
z8ldF9ldANT2lCIPVldXj1kEjAPoXBXs+Yl8740/gGfoKWX+1OKPvb4T2mNChwEiwEGIwn1uEQxK
mXsEjWlTwWIRmULpXvWFaKGi3R+SJk4nvCwXAQfEPOHmiL0KsMSCYpw+VqBobxe2eB143rSHR0TA
u+9mun1stAIYFbFXRn4UpVgfoOx1nmCQ8FRIg76S0o3SuGzN08bI2LT+rpyQbN6zVTv1AHcaJI3O
fTx33JVV4W6bPwwA+7bx7gHm+8prylH5tQaOqIqXEI1FaI6XoDjhaKVeXcan9Lk0ZYyaVyZTYgO6
BOoPUOxfvmETw8U4XCmajrG6oUJjRthBGy39XVoxd+THObsdDTn69zum3jhRER7Oz0u1dSBJ07ZU
ApWGhnB45A2W9E8AKLr1PKrOKjqyAQBThOvTWi++Hk5j5DaIfCkMaSVMoBcJp0lB1M+4n9rtUVVF
mzXLBsINgckN6+mu4mhlUcPang8zcKEiy9kFWnmxVU/cq/m51uQAKFRQRqZ9sKcgJzQAnmF6aXDn
C0YD6b86mAMsnO+4c/lmxUIQS3X510DWWbthZc7FMs1Ex4mBWL4AIHsssEI4dqOk3lghKaD5TMIv
nYsJUz9buTUImD9HnrXsYEl87+y2i1Xx0hVFvAqhMN0xPrqQ5es9jVycFPZKIdvjaqTWfaYOE95z
IxwgOc7CBtnU/+yyzVVAjjtnsZRy1uFTqNOBrfqEm92L43y6IW+zOJeOvdP71DTLq8L8+2XOx5zT
mMtjWIa5kmfhHmak+Km6b7+JgoFJMn6rlOknqs3uNZghmu9Xk77ZKb09XFW3UzZWI6RKXNPdZ4lR
Y2sJDcZHEnF62CYmvIxXcvCkwuXE79sKnfes2yNMY+IBGzYE4sX0jDBqS+Qdm3xgtiBi5WRr8JRk
Whtvy4tOHHuHryqhYd3FFO3Aa4aeidULAYwrnUeCAV/5WkN7Rjs8IX5aWTMmDDi3b8LoH4DMiS5m
VuncbjsxxgLn1a9vHP2V2TIrEka0sbJHcpbyCYgaRHTSh5GGfSm9Dw6OWdas3qyDEKIOx55O04R+
AuwZkwRwR6RQAmXCNarFc9TETc0fm3FnLDAGdKM9qxUZMTpihd8UI91fJgpp0HM5Wghqf3stncu1
EUOnvbupTteW+qGGTTdlrR5RxNFNcPm9ao7UtT9+MsZ7Odbs6J0rjQ7c9ksGbDIZt16p0AJI/qK2
lLlM7/LKdAn5oSZgvqmhWJuZeqfaLUZfNThHrwoHb1kfpkoYi0imGTvYMj9BnJCEWMFFUQcc9fFa
WKqF7Cma7e3ZnkxRS5DWOIHBVadPULhPSdFgIZo4/9rbUW4CXTAehJIXV2x994m7ZAg4iG+ZbUP5
m7+IAj0Svg5WPXWo4QQ2Ps2rsFu+LZ8LfaydTWWe1/FD9Lxk6FJAh3xj1FMUY5x09D4DpWI+SLw+
oszhSroW/kntkDp7MVU3YrCxKIbFFWX0v2fPLU574G3s8eK9JG6Gk5GjLBjhHEpqqFvaeZsaJGr4
k9eYvaNPOhuc2XCVB8unByMALt0Bte7ojsOJMGpW2wRmwbKJ1MqBnnasGyurCeXR//8SUeTCKgp6
dOSiZnas1wNn0uPJJQaBFpSEsfewlOVMbh+DvgkszlX6cVukPBEASs9WTuTeHDnDo8wEHGeMTKKi
ukKhyPnAGpPg6vgcz80Jm7gkZzkCUkxAO+AeI67SW9J142REMMx58+R/LV3om2uFXXcmoUyOxmHh
SicMCNEXsnMiKPL7k4EJZp+yvVPq+GE8NcbA/84JmR82OK8kkermiyoppCZTWT8p5fcPeWm0Me4M
y0W3ZWiGsn19K3bwQy4ejxrC387od8ptho6jVXmWCigWggm1I7EYhuEPDgm4aaGMV8guGF2nQAzx
+yc5T2ypaZBPZOEUXLcJYdfAUVQwURocIgqlyEFARTC0ML1m8oh7bKciuGVGTqhGX2KHEF31J350
ATn9itqHU0uZ0uav8n5VHNt3GGuUmuAm3RT5J3SX9e4la/bjAgWkHV4XTNp+HuNCZ/80JG4DDF22
0hiiyfKpk+BsyoFRCrVWRvcs5z2S0IAGaIEYfcuaEjIRdgusrA0YvZ6Q5L0+KHrNvOAxSz+H2hLa
PJqT+i3LiY0A92hzj4uS4Z/nKGfGIG7VjUOHshSrayZYhPEZ50DL+Y6QN43lW56dGGug7n0LI453
ke0qFf2OBu57N4LCeIVjK7H3KXbbthKfss/RPHfp2Dvbb8kkjbqMDmryqqEr66Ep/02nOdT8dD8y
mMcvMPH11YN2wyO56WbzhXW4spj8NccnNHbIN/QJSTyOE/VAv1g5CwGTKuRjrkCxbWwMXyJOw7Nn
nKbtGLjK+LhR/sQN6H5ZJvUJZSYqXaZfk7ESUd28tboEFX7qCZ5Q24Kyd66RCcCMWAd4DytI0dpR
dmSaX0qnU929x2Vgb7OrPJbXQ3PSNOLMEG86RGUcoU3K5NjzRI2pu1jWVhmmg4MX5uAVQ9mYz3aZ
UgM2EAq9albusxa8XOK8cP0kApPRgoGI+EHBqtWbn98KVme1a6j7TBEhirOi0HLHGtlIT3tdvdqF
Qegh8ZcOXR/njxzVbsT62a9OYMBb/TQe4ymNBg5dHcOltVJSvNFrFSQa3W1nvemNtYoYr3hOz35o
UJ/kx4VyXbNQwo2k9JqkiEcJ40d53KX1U9l9rpBNEMfXrhBZ5rBtgNuS93hpT2Kl3VCOATeOWNaw
CwM929pQxvDyK8K55pHtiWv35czuZGzFBvy4vxf5Qbs6dDAq+YjtC/OqUXBGwj6YqOsjg3DZroSL
DEoBi5EYXhgBjHgCSkivP2EiGYkHP0UoI7o+GvQxG1+wtGQjJUhvUg65/fW1y5KUgTPKDImSYknn
sDCq1v081LsWfe8wsS1EAaeo7Foohq37v/I1MEHi708QczTLAtDKShmiFtho1ctdwbXr9e2mwN05
R5N35vgUhP4F1RgFnXFbfh+M7u3Y2z8y/axspApfyDWApRBiUZf5h3cqXtmRk9l/tBovNkrAURwG
sxVKEcOyh/hQDwUbEgK+4BfuqJAbwgy87OvktbOvuR2flpENLMskHjHFjqrIgHDqY1NwBDNjzagc
g1xMu2dLluCLR7fRmmt9zQ3Lr/oYgqsgo3zYW8pY9Vncwl2wZDx3beuYEpcv8yJ7A1IFB10Qh/IL
qFaVNxy1hyivMtCGQ7mxknSBl/PqsideuM1HgakSUL/gNeIt2RAJJ3y2kllhLKmPeWS2vOgunA+Q
9oDMaPDnyyxdyRe5MYK7m2/EvBxLCWvaVQELyHovV/SbSS2kTaY5GdG0lvQkChDdrg2n04d7azFg
P35ToIEotXybX2HEOWS29Ax0l+BnWj3rD1l35X92iIzQGv2I1rH+zy33QJ3LLdz1poB1s5xvdpN+
g2FfuMaswh2jhSdKC/wV6inCPeAb7pschYNbfhxjncRyzrNt8LKZPeZeHtm41JX1JPHkzIFO5tdV
blU1EHWJtvv05vKg+SFyORnSl5Inle+7hKRQpueXcepuDNBqMdc1EDB3uYwoOFtUNa3Qvb77kB4K
mokO4KU8YTz5Sd3X1Yt5d4/0QzoKbjZp+k6k8SHsKqltgbD0DllnYL0PfPHk2cTMwy6MZWejigNQ
XNqGhzh1lym7manKbDc4Ue26UFZU0kFRd8DW6myj1p4TQt8pmyCKb0DKZn53PUaMJt2G+mfkrbqG
asE9JXH4XeKXJP7mXMOBG6dCRCmpdaEeKYazo2SpZ8tfSurpyNOB3+wHinV7erzUf3IF3BFVG8Df
vtSC54G0egGLC+kkhG4pGrSdQkG+Z6XeRcAR3rlJ03NyGXFMWhxl7QbtQKvzcsc8ocyTDm+C4Hns
y6yLFyXH1yv8WuT76PeS6Ml23mwpqnaS2Ws2A9l2i8OH0K7NGlrVIvTwjkcK3d1FU90mw2R6Zr9N
ioq8DmBJYui+I8a7fj43OSwjBnwtAmTM+8gpFNeHlWJwPL7sNZezmAUMikD5hwVzheDaGweA0En/
ZjzMBw7gP+005kDXaQQencZDAMCsJBgaJrOJDyRPVN5LOOWJSXtSpYynFiqMCSyTby53D7ewHd7X
ny59B/nGoqgm9+xw3s2326wdHxnYV6P2iCpn0oB7t1RJEwIwea2p058zDhKhe5fdJ1G8Y4Iy5CJy
RC98CBaZSyqzbtWaF6n53zf7Ef3hanuyPS6BRCUn67xNbdelNnZQzaPXi0xLEDiJ5CI0+ho/OL4l
E5X1Rdb/ndS2tT/w+mffkn7IVMizuJQAHysAr0FwFMEqmQEjyQX2lUm4c2+DW3VjkfQ0CtYpHMPW
sgkAKmcL2lNam+m2WA/5tdLB87cYVr0DBPb2SvTkEuBgys3V2WmUlrKNtvxSMEZaXIWhC9BxZjNb
E2AKgnmSEtTcyl/TQGwn0B5cs0jMAjvasT96cddiMFko+aypUAw8f97HdcBBNW6YRTqrDYTe1v6A
cRZEwxzdKpcd8GlEz59U/LDIxNXgIuSD/HYbKAsV3xX3++OF0/kkkMYe7spvjv6Tn6aBHv3EV7I9
ZWltuh4LiwvKasiX1+DanrgV4aCZu2zW8rzCo+sjc/JZ0/NtH248iArLcqG/C5nNH/e4rXS3+/gD
Hdt6ioAEKNOWoZZY/1Hlpyj+aFee3yp1Qoyp3wpTkjm/LOjxp4vLMEcUeJ5GxkqGJSFSNZM4Foxg
i0ir3OdYVdY/0dfVNzEzwXyh3u1qShjsA6X0/v21bFGpH9VgplGNT5omNZP7bMNKBWBLvIvq/7LJ
Ct8KNVPayZPmVLjhb8bggj3ue/Wv85LkGkmV2V0vdKOoj+FsRpR2j5oMXxJ2CZ1rF4ufMR1Pdi4D
JhjuefuPuM9rEaHgdPDe1SyEft9SHlYsTBrf/UgfTwl2oMvKhMgAfJEkf4b2Q1Di9udTMWGIV3+J
ftbnTZlpHYaPA5yCpapcP8foZHfRiXR69Ew1XUbrhKvYM0ch0jEvyFFWZTejpmsoOrW72VOT6/cO
pndWZicnf1O0FbSZlrHeiN9ADZO7+njxIvOHGker51sMkyCt+EC2FH/uJtQyx19oMnqJQNhN4oPa
i1o3Mg8XQxLY04nYn56w03RO8Eqqsq6lDqhQT0Jgw8e7NJOtODc9PabODBEKDC2xsYnaFzxvOXMX
uZsdOUXbqy+d2kEKvcJ6X4YxLkflX3VYRX18z9ArCKi/QuFpTyOdUPCBYnVGFyWlVTFZIhNLYT0L
VN0iJKkMHbxP6+BjbYRcbN5uMk9YoW8FrYV1c+hN5Q2S6u3yN9M3BZ7J/y9Fw8vfWtzFzeYF6rpL
64HNx6exntoTkrJb74fqHWqwh/qINMAyKpvhdNciYD4dKiRFYkSZ8HbjlAZ35T+KbVfY9KkoCt6c
0wj1djGREgwZx+RW38Gma93cC9YVX2VdbrJaCEBnBW0McOXBeLWSZWnJIdn9xQ/4im6HhZiT0LGd
ktIVq0XuliP26YgdBqihD6BLoMryEwBe6TlbWqDDwwVQUYnv5yy8537O63SFWVlmu/hDKpRAsmD3
hwNXB5pRV3fNXhzncr5SGcuWzdaKOAtkl2nuErQZXJywZFCD3VMNcAwUbKSJPdmHSIHiCbEQnfr0
Lq0Z/ZVx6kfNv+TRmyV9RxkljDih6LkAdiujfN43g92QrEggaHHNwMw00CxPFG26TiPk+LucToBw
zsxPUZnXthxEfU0KLGaeT9lxvzbUtHQisAVMdWOkYMq1FyXTM5cKcPNNXKnFCiP7gjhVkc2xHOTY
Yb8qAlpd6ovsmMGUUQOxDQdA7vNZTgXMELx1XF8MMYogRWpl4CiqftFk+ltd54b24dJ9guKLce4B
yZm/R/u72l2GNw2Bd8ohqkyoYv3h8bEswkmCSwQ0Be/CGIsVQxQitfJzzhNWHcVStVhs4HC8ghMo
51GoizbCMNiZEjvLvV0w3rgf392oc6woXQBjxDMxRoLv+GnSpOiG7wVW05YQ0FFFrt47bcbfDARq
YrNUD+Tsp/hR0DbvtdJTUQd52wWdqOuTCTJnb0+12UoSvkPc1D/el/3vMcQdCg/DbPr6LBHFGVnw
rpY0cGy69o1QM8vhjIvDj/AWVKayCnHA+4XJaq4fIAlpCI9MMJ7fVzbGFqfcy3AQ5l/j2YitUpfj
+KJUoyl7
`pragma protect end_protected
