`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2025.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method ="sha256"
`pragma protect key_keyowner = "Xilinx", key_method = "rsa", key_keyname = "xilinxt_2025.1-2029.x", key_block
qqEk+Z5ECunGRadhhptsg7aGyUy1CT6YJEBPfbKkWOVZUBjdsK99KfaiTPc/aoE9Fs7VoSLmvTwf
iei72KwvSviYzKpFsfQpvNIC/cv9fXQoW7VRl7kLVzjJMCybRcRhaKso1cB5NLgdxKddHboKqjCb
jg3hu1Ti0DM4idnpTpoE0u/N2FW2J6F1UDh4yVknTnwKsLb6QabjPA/h8RYrkaLoSGW1M3q42L7K
OzdBDHTgMcLHFe9YggvkQV7Cg30ZfNLAmQziZWisp76ouH3anN6aEPSsibAk4auKAMW263HU6tR/
tDtccw/Hbpgloi2+5W1lYw8W20DtR8MG6SLYPw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification   = "false"
`pragma protect control xilinx_enable_probing        = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="1ZdyPR3QG9bk43+4W7fMxwAWVs6bAXccft6wl2DXOWo="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2608)
`pragma protect data_block
Zn0dFHBA05sGuEOzF/ziu/C57q6pJb2NetN0rp9vrQLtcrowCmThskHYUN6lLb73yvrAg7o9Nxng
GZOSY79KibMfCEB8Bcz1Kdsw7JcQuv6JzE0Gvk9ebLaLlSqfWUq2riJIXvguku+3GZS7nLVIG8pd
9kF7BNRuu5hzkN1BgIPmrxFPS28tSeqIB3apzhxE0VWKfJpOqTCDJ9MSObtZuetPZJe94Sq4X6nv
/hOpvpp3JWhvVoG29G5XNaJ3SzpOBjTFzE1VlpTVGhQNDLwnHQnWpp5VV0LNaQ99Mw1n9j/5HxG8
o2zUtBS0uUU/kGuopAJFcgnqdtrUqpWiB8AtOirPRR/vLgnjO/Prq9miWxRRiT0Pqe854jsEsIKV
NYRx/5z9HHlvmBFk9H98+UjaBZxK/A6x2GB/GOgv2wFPDrSANKb0Wg0ay39U+3A7GGiQ4UTTPCHv
wPcIhg0bFrIg6rfyVR1sMoHSpKJP55qvQ7QJWpT/ifXO0OQZ0jRR897+B8TkLVN20i5xRdtvUqUt
VSELj8uEM/XwNucgt3jTwDHUrCBAdv2sJqR9lKotFxYsh5KaO2cXTI3Bspws+HTgowCRPkbXIQC8
TFRhDEEiOU2euP3QrArvbT1ceJLOncgiv4g65tE2jUNUI4nTBs+oD/sa2N0d/Uzu0CE0SOktX1ML
KUzITJXQx4E1+bHbtVmGcS5KT6bwAXBCCT2Y/jq19/mUgOnwKUkH4V2uRfaC1GWLI6BIJbu0XXEW
t0nMWf1nlR+5T8AyyFiLTn1LvAVFtJhW4jLM9Qf3bL9ToTjPtLb+QNEdtBhqq2ns+DplbVmhT9Iq
l3kDIzybpghybtFgDJPckdGuBOWCVJKsEeIATozC4NM8NYqVnK2wlkvBowuUPlvxch+VtRnAge2D
uKiQmRSF5sbbNZL5P9GRPRfgB1wO4CML3YSEQiyKbPhvmkYYfEGkBQnMuGTY5NczCBoLULPybMfO
DSAKF+0JNw3BrgFX9EYMpQ5lcR3obHy+I/BBHUG8tJnPufEyEKiPcgQ8dpHrAkOva3EjH5Q9DcA7
OeFfUymWALR3Lgmh1YBTJWxBU59ufcDP6y0mxcpzuj3vVtpipu1/U6XhnkUwLXEPRKqQgd8GpDFZ
j/AvKC5n/+8C0w7+hg5nFnuHux5ww/CmOUOhLnaITmq+FGDn+N5iQIht6MJ2V6/Nz76CqSjYG7Z5
Gol/mbEnomlr7zPmyqeRlMzPdYBpDMwx4ATyrgH7aYqygJJb9yMwueozJaR8ciIdH0/unwrpcI1z
UrU7J1Yy3fC9JbgM5qepIDMYwE0LWrZh0ro8Wbc2AHvkmtQJUrRzcGmIogaBIvuQZMHzLbv47IBh
IJg2Zbpi9jMXg+zQNR3yPptWnPF/+Fgr/VrOfyojNcJJkXIEBRp6+hCR3OTiHT8e3cM75oRUsbBM
Wjs+o4o+VwhKzr1T3ap1Q8xZSmNDNYnjKi6PoZRCtGxQVzG+03DG7mGKLkzjjOdl9Xo1F0QUpRCf
f0zU0FzJ6rl8xWJJOZBiq8JlxVVnd7Nmu/+eW4uNPqaenqbwCPxHC5kjZUdHsTRS0P40GolxWP9E
DJURJSQsm+zWR2PWclhlv4SwutKz/VDEF5zk3bZzdnA/v+FHcN6STWNiHMc34tFHXgfb+zOWeNDY
7R6pQjczUwoQEoRyST+QO97OveoUwT7PZ6bXX9m+PBr1uuKM733Dlk808zWTHLk091V8x2x7XEq+
H7EWl3YNWPy74BLRwjJdwpf+ManYsir4Vcy30L8ZJS58QlNLw8TgJxuFT9yZ5dpZPHt0altZcQff
zMlqJykO319AKeLkivGBrM0ngn3qvYZI0HGoiCtq4m06QPz0Oj7MNF/wqWdVAYCn5H2Ga//8Tts7
RUagzE18m8qYItoh7YHVKgrdhJAuB1nnRXJgNp8nSV/L9VytS6XR+hR52RbL5yRSOWJJZZo5rnsd
7qTdKPaAbrSwFYgQLfTP3wSg4kl3X2+bEF0fibfxZsUJnS6yugEh+5+72wHn6e6s7gIdMUymr0dT
okhrXWn+9rudPFOh5ZTUhZ8JaptDEMzvBB5aoh8PNklhuMD48081ZYahIRAfZCBWf/BM4qOZhITv
BRjAWJaNIZyOj8w1+xctgGqgUuYYooppWMicKDGcWymwzzgU9oiLFtzpMCgMff5BvPgpe12UIp7J
2KlFREe8K4jx5Q1csYnd12QnaO7qqnHKTzVodB983NylH0L/nceI1aqMmW+u84Dt4eiOzJohJP1a
3Yl+Y5Wh4ZhklpvnKD9ejvkagAU81HH/F4ieMMkzV6hxs+FmnFehnnhaGWV0/QVwFrdtWwp7glG+
Zzp+kWw6QWBpnfkdhxOHJMghetelpQO5oNIH0rdPDb729jTm4Fo/8jcwmieLcRjJ8fzKepQuf8ov
N2EBWGz3JiieuCA0Wm1Ve8Lamad4DSH4VQJiAOOE6CKjAZ06flfd/uH0oHa/QSmIRujkae6Gzgo/
4s8tC6BcaUIOkLLiHAHA6pk4oLgrL/xHE9v0x+Suk8MWEHVbhbOfO3nM416MClKfVSgg4vJy+Msb
CPBgPUdw8wDSA111RHP7HR577Q+MwBqsei6dbckzqFYjMbi6yZB5diZg8nyfGQ6EQdrWy/xk0rb/
rXhu5hw2FkhxJ6JRwMVloEfyJlNe8kbA9xmdJ7fa9xj6lYd195S/YleNJVmxeVdHISNTPXc7sHJF
ZsHM/3PKzEepa7FjsyCWPTwUw6em8aENdv7JtgOTeinidzd/hvF9TxaYpO8jFuhePqEkKX6OAnNQ
d1xeUKuZJqQxPHW03AybDMUn0FmQ1HYAqJoJgVJoWRNo1lJ4VbMkR5XXkzztLZUAkg5BO5+JfqBi
sRwAqAI9ZxccvmQqx6YMwLRUlic4BjohkgeIteDdiqdzbvatjpRVLX7CCp8WRjmSsz79MlbdwDD7
eVU+Uegzf23iPfdc9ws0RVe2S08j9l5PCoXph612PS1a4mh+2Nc2GZUiNtsKmmVSyVOtncK57Znj
HvYJu1pH+vz6a0tfAweYCqFzEdmOju/2293J1l9LbWWRz/vyhcVYQrp6ufR3rP05o7BtmwVOv0MR
5xgVKYMZGw6B9NOQm1bCwziCUfuRP/ARUmEB7Do7MszHLv0htwdtai18abeQ/SZmF70FLiBa2wC9
4qfMC6AkatTLbPlRV16nASMVmODuimiYXY/XF5QLEn+0mMpxaqFTnLskKjRBlKDKq4b9mshCEq+F
6m2vnQdoYm+8uzB6gOt9E9p24jMPP6k0rQ0XfxCoeFXs36v2vKe3dBbo9UCSPkMvqmwD8LswsbBl
oyUUnMdj2809DeQ+aUMVmfBUQ37HBIP7RP0l7MvlG87RfDdt9s6vSVG5p7lxx3aa4Xu9DXRg1mvg
2RoIDrn5Zucbus6XBErCCBu103G7QpQWiSKndxUiMZCeKmpvm42dFq/85A==
`pragma protect end_protected
